PK
     !F�V               new/PK    ���Ve��2�6 �o=   new/SETUP.exe�y@V���PTR"L2*���:$"���h95j��&�R�Z�#��6hzͲl�Ms@��Bͺ\C%Q�n�0�f]��>����F�}�����k��g�׼�Z{�����u'��_S�8[������1�7������Ϯ����k��8%j�)M��<yJj��c���M�zxrT����G�<8��ƍF�aJt�����zP�w��mP����|hg0��8����PE,^���~���J �4�gnǛ[Q���*]Bm":�\b��@���@畛�ߜ@�:��w:ʌ������/��ߍ�cg����m���������/�>s�����^l��h��9��i��� �`pr��	��_��c��3�Hgy�i�qe��A��SR��#4:�o�;��2oD=�S��m~��o2Խ�q�+2u���_�$�u�p���]����L{�qDfs��F�Q����<��s\ݸ����~�8���+���������YѢc޸��\�QXof|�UXo�w��J��5�5��~��v-9��*u�k�˪��������h��eQm̯��/_���VVh����y�!��Qf�.axj��y��Z��1cݩʾ5=�w��	�1n��F���?uҖdn�����|�E��EǼ��C��;�^SS���c���.�)��t����%43=�I�SCM'_V������gIj+��WM5�&D������V��%���yBt���r{FG�?e�l3w�7�g�����dǼ�G����9|Xv�꤬C��^�"Q1���K�~g�����.=���&��$Np|3;��_=
C�E�q�ʌ�9�Y�Ur2d}��p9�تI�ci�逐y���|��2/�V/�/4��t�|�_2��۹2
Y�p�r�w)��0����(�"�lvs�b❚��C��k��N�����FTY�|A��U��0�̎{|.�����?5!����[]d2�B6��95���O3�0��!	����sL�p�!����c=����|�U�Xij��ݝJ,
����z͉�w|qe��ɵ���貱�羫\9e�~?�`�^��Iր���˲�f%.�O��I`fA`��ws�#�g� �5 �n����Κ��?�߆9N��K�������-d��j��U����r5���Aó�:Fc�VE���r�t�L0|�5v���=!�N��4u%gtz�R�#cO�=r�=���.@/Br�O4�]i�6xkd<�귚#�Hׄ�G[ҟ_缹c��W�g����v%�v���5㟾�U�_��q9Y��5Mۈ�O�͛�l��E�Fq\���kT�L�N��81�@��yb�A��A\���
�-��?����&G>��N�r?�K��r������s����$�˥��xM���Q����5ֵ�^Q~�n#x����"��PfEP�'nK[��@�e�O�^��h/f��@;h.�45�?���J�~�CL���U��
���Y�
Hy��(��Um�y�j��^{
r��K�%��lv$��)(��7 ܗ��m��o��9�fA��=2�0��ɻ&���^���&Vr#(3�: 3�2`nF�����)3��p�u��gfT;���j K�[�Nd�1�K,q%*�j�Z�ުgn�Jp�%�$khttv��'��j�w?����7��9���sS������T�����Km�e�a��Eo��'�/�HVbEab�>�#&.�^��'Ԟ%����c�	�I��ch�q��9"��"�׮��W7��%�t���ڲܝ�3/,tz^5�� ɗ\�=/t��^v}���u�{'���ю�3��d
�"�\0�2w��\���K��c�:����Dw�q�P�ZPK>����s�=��X�/�2�(�x� �n�N���q/+����7$�7��ww���e��������\j�R�[���,u�Y�B�Ι�ug=]�8�����ū��;���nS��e��a���¹;���9���%�j��y.T��=���1��&۬�7�U]C��A��'����\��O�L�H���
CME�Y?�ff>⶝46z��k�{=x����>��o�m�o�L�Z�˹������J��1��BCW��֠�A���.ԦӣS����z?�J��AU�\8���Sˮ��A;/4�iS�N���A�r��A�t�]ze|�Բ�:躋�^if��O�+��A�4�k����� \*Qi��s�"~u��.vl��pjT�F���?�?����? �\�8h���lq���zX���&�Ӣ��;�B�T��"
���&A�W��Y�$2�Ĩ�k�9�-��Ꚛ��J��Mk`��928�?�Ukp�;�]��r�Ӧj�auz���z�W�S���]V��n'י���N��:[�����U�,O:���������~��^eE���A�w*r;�^��t�>'�vY��q;����SU���Ǵћ7�۸�_a����3(���wu
E�V�:�%f��9+uUW�+�E�p�D!�q���^/��:(�ꚻ�j�^�y��0�[�Va�q�sĹ- ��%���D�E��ܗX�����
%�ˀ�&H)2����ܞ�ua�>�`���%h,����.�l.�%���c�Veg����//;<�,L�#��"��i۝Yɻ� ���]@n�n��i0|w��&��07c(�.D)��sb��$��t�$��̀��d������ ����$~���^=�Ƃ���<�Vp�S���p���CWzy&zꙘ�\�7O,�[�+���͔f���(s��u��{$9@�?f��rR�gf;iC�R>ʬ�Y�վ����x�6U�lv�/�\��*���L-�;i����2M a.��-�_��}2���`p���k�ئ]*mf�|NZ�{?de���"e\х��T���T����F�n���^~:�~�1ӺJ����}�T/�v��y��Q3�6��� 3�#�&zuR[�����L�n�\U�&�
��q���ϋ�t���3.��+�a���4�tr�(V���J�z�+��PC���G�{�������|������`�ăLǐ�"�#$גt���E�����a|�C �G����B�g]���"�:Ft�B�����"��/��"��߹n�_@���h�@;������	�"˛�}�q����������g�X��l����5�1{`�����=�?w�w�Ѯ��&�����Z_�ia�fcn�Y|(��e����JN�L�y0'�7Z��i��������x:k�?A	�H�XA�w=���ɧ{�Y��ӗ�� G�����ϡ��C���迹���,p5�_r����ՂA����,ҿDh��������<=*�ը̼ m������o ^<�h����!�G]�5rx$( ���f��J�5utmC	u�4_�2�� �A�~W�>��ì�1��>�3	$+db����K����xܬg��#�*O,Cy+��&�01�/�MV�YY�]f]�U�E��u4	�)V%q��]�3+ߺ���X�쐱�,�Û�_�����$�&���Xa¢�+3��E����x<d��B�X�'��_�`W%��4��c�(�2�H@�����Z�?}˧(���|��:�j;{�/�(�J��貦 ,�G��Q�x�L �Q]"*n$�#����q!��9�\�")</���笊
Kp�bqjKc��rj�h���j�^�>6sW��?/ܿ0"�wUh�x'�\Mj�����ү&|��i�&j�io��rc�"Fd?�t̓�\V��_�|����i'�?�=���.��_�+����>Y>ϭ7v�+ȱ�I}2:�t�T7�	ũf�j�3X����74�EL��`������~2����2�3{�>�q�6,��*�uR�e�H�#sW8 F��y���7�����q,����u_]�U�a{K����f�6�?v�M��2�qjw��?,i[�5n�r�y�/({pM��z��Z<����h|�oj��Q�}�Ƈ�?�G���E�S��MBz4!�OVjtp�(Y��IpoF��x����0����вzM\��v�9F�(�Gm|\��O�=*:�l�d�AW
}�J�[P4��mo�8�c����\D��n��l�i+���ӏ�Ò�
U�����*ʩ�g�e�%��̞̼`_h�/�5���;<��!Of�r�0���i�d��.{���
ݍ�*�?2�����	(ɚ�.�fƏ��IS�^�ۃ��g�gGJ�b���Q6va�Yf����T�Ug~s.-4���g@殘�c�)�ct�7��}���Bv���^�N��/(+)�������p��3���i�j�F�V��Z��({漷I��٩͌K�,_Bp|��2���v]�(���"��;�q^=����B��5����������� 3c������p�����h��l������2��|��g˽m��_���z��T.�<��6��k.!�]u���^^�e[*�ufA��snϐ��Y��n}O��e?�VC6��,-�����O�9�o��	���Շ�QiӍOl{�.��~}ܕ�'!�u���B<�JS�C���(���27�4L���0-�ݚ1��?d�TW48m�����j�x���A�:��ݧ�}ѳA!���� u�V{ɵP2abz������'}i���ߓ1��3��&d�(s�y�LI�s�XŊʎ@�r]�3���nr����4Gv��m�6\�jUvڷ��({v�GفO�B��Om�K0�7H�����n�Yг�k�O7TB6[�����e�����8�����K��Pv��\��q5���N�{�N��v���0­�d�OS}=3���p�g?�i�[��AFL�җQ|�B|W
G\;���]��^�O�)�����2<�˽�J��XIB��s��\��J�����GK��2w�^����;��ǃ�r*멁��sz����^5}d���Eȼ/\F=���]/���w����-�:������y����K]���k��3���5�]��Zb@�=z!�^&�C�?s��}"�w�{�s�������[ƧNugͨaS����ÐW�\���_SSc�u������ᎽY����9��;u~?^5E[ܭ��o,|A$� +����c���.���i-�yƀy�[�����w�"�`w����Y���wC�2]7���Z����'5����*5�8��.F|#�旦�zк�>��;�jsV�)����e��.���'�vN}7n2Zx�A]7.ɺ5���\�Ѭ[�j��1�YM(��������:8�Jh�1���Z�s�$��ۺ��F��||��b{6�"��{R��L�5�皚����/���0ˋjŗtuB�1-�o0���gSȼ�Ąo�� K"$_����N=^v����/->O��U��{�����7�?=YScd�Sa���EL�s�y��7�gz~��ߧjj.Bg\N�;�7�?�}�@t�p	+~r�C����v0"�Q��ع��s?�AYE����fD4
Y��4�3��C�Fx�u�Ć���;�~vB��qF�w��l�u�hhZ0�P	���]}�X�F�3�c�����A��{���F_t�I�*-q��"�E����Br��Ko���٣B��?�v�x��a�'�mz���ʍ�(P̌t�0���{��CV�`�OK���a��_c���᱈�P�<��3n�V?J?ɝ������������rw���?��a�!5��wT��>�N�!�^t�K������
 �<"�"ꏄ�qs������),}�+2-M���~�ߩ��Q�����<����H;a����?ğF�^�^u����f���Ü��`W7U������������2>$�Q���#;�q����0?�?7�ߟU��&�9�j��YE�c�p�a.�Ћ�"�Km<2k��{<�<��|s�8�9�;��ˬ��C/7��I���)��=v|�2�\��٦G��g��1Y��)���.��5	of^��O��mb�7,�_:���'����|b�ݿ�H��r��f����t�	�:���/7����7w�m�n�*1���o�?<]�F�_��W�ނ�4մ��\����N��������;��w�����y���s����������������o�������Z��]��r������5�?ܿ�q�8���m�8a���8�r�āe�ng<=�9N��-�q�3,t��1�b�{(Ϲ��F��rk#ÍC��q�s3���q�p"z��:����0�v�Ҍ��d��n�\4��d׆>��E
8M��qZ�%��O8�@ǹ�qL���qJ�����j(ڋ������>�q2���D:�%���tg"Ù���/�d�����M~�4�i����� 87���m��N(w�:���Lp������$@���,<ؿs�q���)����8�Ha@&���W���,5���<
>q�S�'�;N0��8S����� 1w�W�CL.����8�"�L�������>+��|
W� ]����ޡ�1�y��; e�^���0���� �!�����H�2��@�0Y�P �r�Z������Wi\�"���6�����l�?�8?8�~��D1�.ҿ� NB��s8B�íW���Ĳ�0o��v4�QH8�����T���!����p?� $�y���`:j&(�~a��(��v����K`2���c�.�Ɠo a��6���E?���N1���\gѢ������p?A�#�nU~s�h�ؓ8�Qi�~?J�y���Z��o@u[>vg�����O` �0s�9��d�;1� :�2���߀�E{�y�n��M�ꣀ>%�Uh�- ։[�P�B���zPa�Oí�t�=*��߉�{ �0�� |3�<�
Lj>ζ�^�ۓȽ��U4�.�	��x~��ip*��ގ�0�p�N0��碁r�&��G>�>��7�����y;S� jD݆}=�+�@�@N�I^�F����N�� d��bV2�~��ea����
�o�	|��J��e�zػH�Q� ��g����`�0�7d�����I�3�y;��C]8��@wS���M��9@�S�x����܉��gw�	daQ����M:�п���V��(�A')����2Fu�}`S�4�����n��_�H�a�-�� �H����@�5P͹;�;�]7�]�T[:�A�h�o�} �nQ��@1���䑪�q�g5�>q��r@~ ��Jo
�_�wg����@`��� �N�[t���A~~��M�B;	� �I��-=It-���>L�F0����$��������Љ����w�K��Us:�v�(��*�0�u��L28?��u3NIAo*p�3�t�R��7J7r7��]�:�q:�#�,܈��}	4�p���P-�-ѥ$V�Ů��Pe����$��^Sٽ������G���j�/�͚���6zкC�H80���+��9�����F��e��{�9�&��Hxہ�1x���qJ�[��q���o����}F�Ō:L5	/7hf��q�������~�����.����?HT`�����&��;�h+�C���Xw6YɃ�H�=�@���8߳\����Ɗրu|��u��R��W���Hx ��a�f���V�l΂�#.����ώ�Gd���6��֠�>/��H�.̂���)T���hp�ȲD�!���,_�����tb��D���C+"���0�Jma���$5�����:BW
�(D@��6|��Md�c��Obؑ[��c>����"+��!���3&"��p�z���Ԧ���	8M��q�g`}D�J�1���#�Hx��<N���`����/��%)x��n��k�]���L}%L;Z�6>9�d�#��U�<;`�X�B�-DeI4��̃��m��s����h�O]�Jc%:s$����Ё����e��T϶^��b|D��I�@:?��t�ڀ4� U)����0�f���nέ�\J%�hjSϟ!-=�[!!�tr��W����S`��ꚾAdgѱY��"fkؕ�noBg�4�k���W��]�&	V�&�|���q���^�#u�s!y��_O�'�p�F��?xҌx����$����}8���2F=��O�	7b������у��D�4�d��O���Vӳ��ϐ���2s)�;����aq��~�����)F�A>;������Ʀ0�1h����N�\�Ù�u�-?����a�\\� ?��AT��h�|�wl��uД'���4|��Ky�=�[I�?�B�-h���>��]�7�3������i��]$h��\������!�(C�g������b0/��{,��%�ɷY���������Al`�b��I�'z?����}_��v��{aQ'譏�n�r��P�� ܈+W#,*œ������>�9����`_���Ƭ�f���z��-C�ȥp/�_O2��H�0�O��p��ۛ�t�O
��Mdҍ�q�6� �.�^�[�~n��g�����0'�~�
�?���po��ܒw�>�`Q;��/7�� �Շ��iz�y�4L�-��p�iI�N����o"�
~K�G]��5&y��@�U�/g:Q��x���HNF�%���B�cH��d�B��(�)��%��u4z섔���N�y
_�2S��@��1>����ߒ��l@:��@YO"�m��e��1�&�f���n�EaJ2�pKԚ�Ģ�qԑ���Aϕ`;G'����	n矰��
�����70ѥS8�DA��$(I�E:��Y�x�����.�)2��,hK!+�=�N>����5,Ra�[Wå'�ŉ�\͵��P�2�ӭ��EX*��(R����C�JM�R�m�`8� �[��d�`!�$=����n|���W�|e`>F�A�y�j��H����c^&"����1�5��nBp���N�s�M��l��|V�"���p~�x��bc!�jM�7����,l%Xm�-qPT ���n����$H莸�KKAu��Ȍa�]��"�8���p����=���o��-�,�gVba��nF-3H�$�y�w�
*��ǨЊR�RI��f3��t~e�X�J���N^���ؠC���B�|�Ɵ�^Ig�C���
�Z���Y����Z��]�Q�+�xZ�%&Ia��+�X�_z����
�\M�x���n=��=����^aD�q�K����=Yg�����U}����r&Z�t~��~:��Z_�����p M8�+�^�_�_-e�ۣ�_�s
F��p�@���X��
I��-c`���(@<��/��qGOrQ�>��W=9��۟�}uF.��HaN2��fk�9�
$h��@�3&����g� ��Au&�_$���q��Z_����2���M@L4�ƍ��m�:,@���J$8	��0���?��me��ϡ���>\Vg`vaH	��r��$���h��N???�сB��ֻ$rɯ��%��0��tA@K�[,�`�B��i9k8�
��H-Ikk�H��sӒ���@�ì ����$��рMg��KX��C�[���7sQ�� 9���j���T�.d�s$��$0��V���g�r
�~u@����#�`S�@�
�ÙHJ���bC��]��Y¸(Q5~[���K2]��T���,@�0�l<��@������}S@VWв�&���h?:_-R���\���b��!����p�V&�	�S������+��ά�K��,��
��P���6	�ށ��գh��wcH8+HK��
_ԛ�P�#��
�,ƘH��� ��S���߁�+��$ԼT��,�L�ER]yD3��4�L�+�'q��"X!X}�2�	��p!^�jޘū�K�}a�Y����Wu���ux�:��D�9��b;~�:�
�s����c[Ѣ��ćpc(ݏڿ�&��!;��	f0l���u����0{�gQkG�S-��-w1ש��u�ZTD�O �}��@3��yql�ݰ��0�7���xZـB4��ug���0*�Q�j�?��^��}s8����j�*�b��J���kT�a`���Ϙyc`.B��a]#����aI�-�Y���"u�kX�~a9��h;>j<�e���[e�H��_0M
D-��2k�6�A�CЄ��]��K���"��L���C�ۂ���jQ�%�HL�(~�*�_J<��2�#�>������uC��/�s+̔,r��D�Bu/f<�n�OZ݈��$S�Ǯ?�h<X	r�
���F#qɦ�v��!�e���6�A�����O���W�s/<Ïb4������,\n.l
��(�[L�Ӹ����c�B�[$8�񧔝��X<�y���C\g�0�1����G�.�/��W�6#eH7l<�3��vB2�V��,����ܮ�X����R�U7g�q2d2����d�,�)&*ocq\ף�u���3DV�a 6�eH	6���NE�
��!�(blS�@L�'�|7Hc�t8&k�J݁���n�~��R��G�,+a� ��Iv�z1�'ӧ ��,C^�!�В�2�R8���������IUĦ�0\*�Чꐞ����Ðf���fH,+ړ�tgK�!\�AF�m1��K8��=<�Y�aA=q�q�K+#���!�pncu����+Nr��g�끄����,�7a�2Y�e=���3K ~
����5�z+���[h����C1�,�[q���D�X:��J4� ��A�phi̐ւ��	�w��pE49�n�qh�0A�-�xCB|�h9-`���	b�0Dr� �	bC�^b͘kF$��4��r�u�$�r��4���_�^ڃ�h�p��
-�k.�4.��}9R5SE�4��G܅ȥ5!��*��0p�Ғ��i��lH�f a�o��5��u����ۆ\ځ���)�a^A�9kS'f�e�=:����ܣ�t�[Y.�q�﫺Ͼ��(C���~���Y��5���c3�-��vf>�%k��EW L�Hp�����E@l,h�f}��{��t�>�7ѵ����v�g��8C�v�GU�R�R;�LsHFñ&i-�&=B�6�����S�b�8��c2�~�X�|'ˍ V�UvE��ꁓbr�D��Z;�Ţ�&t�Q�QВΐ��d�a*���~�3�h*�)���aB� ���@�J8?�*���0d#r��ҏS&ˆ{G��領��]�j|�I����� ���8L��0��e4��˺�25���dH
3[+^��;�t�e/�A�=-�3�Q�r�PG�	�?S�� �]�h�l����z:Ȑ��m�d���6��E�&���RE�!�H19.�}}���{W��M��D,Ri��3�]V����!�=�QǪ�����m@�8��*������oD-e����e��X��"Q�y5\��	�n�B�!�o�B�P�s�]���
s��J[O^�^	-b�����_�yS�z�i��Y���^����1�M�ÿb�A�C�<��:�M����T��af��ZD��TQ���8G��a�h"�5�ꤥW1�� ?�LWo9ZO���,Βh�W[O�_mj�2�ZU�b�����F��:����=vqJ"��L!��Ydq6p�#9�W�?��'@����1QQ��z�,����AL�*Ҟ8j6p�C�5�\�(gXn\P�����/ݩL.`E�
��uy�"0��+P��Pљߗc���c�)T��YW�U��c��z��"U9�(Gh~%�Ӵ=��h8z�H��L]O.?����Z�y�2�M=;����j#�~�Z�F��s�c�f8�*�xÁ�]�B�yĔJ���ÏmT�� z�+�]jȱ��$J><�|9�2��Bf���*�+�[>b����U�dce9
��3p}m��I�P�Q��,+�0F	b�;�U��N��_Z`�4�iȐr��W��)H�4a����&KR5y��%`���Y����!�t��	�r�� �3���0�Y�ݡ�ejb��,���򿡈mԽ���k���[���v��^�m#���Y�e��/��vĐW@�h�C��a� +jY��Ɗa�NGk8*�����4�$�Zsf��S��<��=���X]��t���,I�E� rX%�"�,er
��yr� u}U�2��.��d���A�;@+$��,�`�Έ��o����uShEg9 /�_��x����,��1K$��@uO�O�!�Q�v*�bp�9����.�@~W�~s���-4D<3=�&�r@���"�\��^�&x�[�0�R�0�q���V�Ù���'T;	�(�d|�0����p��x|��k� �Fth����W��S���r��&��b�*-�0y�jr�,�:_QZJ2L��V�譤e��H��d��(���*�f��X�L�F1�Ru��%�ԞR�Ip%WC]��ɤ��(��KQ�Z�h��$єx�}�K�ו$�VU�zf��,ŚYL�g�:0K�.�^&A���)Z9\!&����W�q�`j)�`-�<OfW�~���ϐ��ɗ�ʼ��^�@O���Cp�]�\K�^��o�{L��P��&�I��6�Q���>����<�0�+�oĦ���,d��C���΁Ixe��y>�%G�	C~%��X(��D��B��cW�7&���v8�����"�
Hn��"[������&�f�nk��;A,	���<�,�J�C.)��R-J&
���w�HB���5ZQl,�o�& �h�1���w�U$��C$K���c+x�r�&#��c��g�/�t���1�(�@~OF]b��r�tF�ʡ}$�t���p�2Fxق��o�fB~�,A�P��Y'N"2�
���
�����v�ַk�D�8���=�:�Z�x#5��Y���UC>H��1yճxL,��ո�͒�R�bOj,ǮDa���бG`�a��R�9R�8�r9	b/�n�ҍ���TȿIO�]ϐ�z��fU���"1̕ZNO ��x��P煣�jY�0�������V���@E��K*E5�"[R�G�L�O�5XO�Γ^�B.b��4��Ő%�KF�i�Ot�'��0C�P�ĮҚ�Af���
�Ecu�
��#X��5�b�-V��+х�����ty��.���^���n�U.gpӉ�w�\�P:3��eC$)��ͨ*Dk�� ��Y�߯��l%?=iD�֌�w*�Xe�Kbb"�fX������&:��P�_V=�RD'�E�R�ۑk��'i*�m#zK�a��8���
\�4��^hݟY�$��rL����n�в�eW��b������?͢�;޵"K��b�n���xv��p,�J�@����K���=*u�@wQ	�hH�<����eE�@c��H��&~'���,�LL*�Q���б��������yCb��нWq���� >�޲R��J�����C^���E�:KT1Q��:CJ��ݔ|�؃�2�Y�A��:��XV��y������H�+k��� ��AJ�-�c+Yėi�"���1��U.BKgD/�*��y�� ]��u�H��]CYF6R�ԙ0��y[ώ5K��R��c�R��쀽��!±�J�7KX�V�c�G4�+p����p,����K:�I��e�f�*"�R���'�ҵy�4�v����Z]/��zl|�V{�)�f��8��m%�T�&y�����L&+�k�W��I�8V�o���g�t�~(�"r�q�K����W�6�3���ų���G�jG��)dc�*�zJj	(��ڳKw�R��+�&���=`�Teî���]��Ľ+�t���K���5��Uv(:2�ox��h]���l��b��]ⓟb���EB뻘E��'��C,�1V��hQ�Z��
~_�fu��doc���e+�=�-����$Ɉ��د��K��[���J�9L�es�p��Y�JF2�
��Ovy�Ӑ����<�WR�kƖq�:%��6��K��y��Ȋ|���P�N�4A���e�,�O@H���)ʿC��f�1I�$��my~q�b�(|�Hq�+C�Zke>�c ��l�$�=�d
��]I�PE�0Cn��'X�&3��m��u��5�=� %��T�gH�5�
� �F�)�	<�,�?�nӘ��Ӟ���M��Ch)�J��⹋�0�a���n��t��G��Z�n���=b=�%i���F<zp��o�� �Lɑ��+�^60�.�m�~*���i����(-�I#�js�Aŝ�Ib�-cu�o�O�J�҉Zq�n(,�������`�Ԑc�|�2y��-�6~D���V*:�Yd_".	���!��'��T��sN)D�%� �<�����Y[6���$�I����A��w!�6�,�`�3�NK�]���BK$��zHf��N�!g�:������z�G����H�sF�]���'N�H�hR.�U��lb6�
I����0��VtI����s�զ����ZJ�>.�I�l��fOWu3����y�Da/W[޲'�ĩ�\	�# X�C������|�E|-&Z'��󯣏U
u0L�+n����]T��$�ʟP6q}���9V�_8&��X�R���RØ%Bݸ��G�0�YD$?cS�/V�9��
w�ک$�q�]+ǁdy��V)Ѹ���5N^D��Ug�Gz�,� �K�j|��'%j��|9�۳�q�UD�-U��LTZ�i�7�YD���[�_���S��j�])ڷT�
�TS��B=�3V�|9�DF��o)�<�"�<�����"
SA�����)�S�Z#@��u�Z"LmE�� �O��"��0P2�_99E��2M��*Ǆ��.����"�L� i�N��\n�ef+%�s:���OR�
����ېG��c�4��'{C�&6SZv���tE�Y�����k��ݸL�
e���=QC�w���l��m��7��Ġ�"�W9�镠�5�\C���::+Ͼ����0��;RuE���I�����kֳH�X�ɉ�����巘m,�~M��tE��-�|���|�00;��/�%i�.�(���~c�4���N�@����S���'0�T�M�'�g(��8y!*�COW����F< C
� �e~�&�_�rZ�C�*b2����\+$�adȂڳ��@a�Jj�t�2�F��"�E瑚��rH�2Rg�da���Yb�c]Y.����E��V��T�~C����`�V�[6bM�Q[J��ڪ[���ˉ_9��G�% �iz:�Ms19x u� �\�CD�>'�ܪٙ�b-��hٯ|]��b�b
Iy������@5�Y�\%�΃��N�)V�R��zpK�=K��jI�9xЌè��H���Y^�Y�uX��"'����S�-�#rZ�;�?�}u�,��� t��	�+_1c=��΂��G��t}9��H�mm��J��;Z#���c��E��ݬ�rNt�&})k=�]L�X�y�[���zf���W\o�[�����s���)�?��{�m�XU�H��LbxK��W�c���ԍ��ॠZE������R-�z�<�Y�e�Bʿ����,��d�3�!1l�}�]��Dk��=�b�K����q��R�V%�!w��p,���eb���]�� ��Dy���֐�(�r"ό���<Ċ1�\� ��][.�1�$E�g�Ej71d��P��fɃc^<�Wn��R5>��S�,���,^R���@k���-��9a"��	���ֺ_E9�C����0/aȯ��'���.Ϸ�1Tbɥ�!��a���kH�V1��L�W3�*�˵B�C"�B"�?
�t̥����j�R�Ǌ	��-�O���"�@�j�k,ZV�^�D)K�a��1D���?�3�!�XIm�� 1O�_(-�X�c�5΀��d39ޚ���F}�]�Lި�L�3�TZ������Ս�1œ�U-u���.="1�U����h+N�QoY���A��Y��a�������R��%}J|%�5���,wq���nqJut�β4~�Z��e�ΒĐ��e�"Vd��m���u���$�ێ3���w��E����X�W�t�4�x�쀖t��w1�ҍ��X����<jY�ܓY��Z�ZNgeW�E�\�E�NS�X�p,�!��_I��X�V1�8���,A�Vk��T�_��B�DO�WZ���Ҧ�,��0�H�������:P�ɍ��5��dyÆ8XO�r�]6�����ݴ�7���A�xL��"&'T��Z�ڈ��d!_B�!�s��Z ���.� C열oT��s��U��9�h��r	��!���C��9�ў��l��=�3���R��gyE�-+u)�e�M~���7�a*���� �Q���#�v��)��4U�GQC�!��eC�f����;w1�v�u,��C��;�f+-/�Z)C������z��M1!?Eg�h����CBk�?՚%E���e�ڈ���/��$}^L�8��$��X�?�
3��,�@�L��Z�=���!r>��!^��U��;�)�HF�I��!U�����UZ���8��X�t���� �\19�9G��p��6Ƕ�!����2���0UE���:�T��!�c��x]R��o�c�3u	�0X"�}��b�&X��J9y�CD�Ǡ���-�������{r��]u�Y��u������VJ.�,�����im|�$� �h�/��E�*L�n�MӀ�Mv�E�+��9�u )G��P�����w*ɞ��a�^��QLg�e|�= �D)���j�<�#;��k�d9=��M^�?�#��� �"��F+�d#���m;C~�>/�Q�,'*#-�|�Y�Z���,���Yxg�G#�v-�ț�� ��> C$���˛�����5Puщ�EL��5D��r�?]���P��M�:�y���,/�����@�np{�����"��$�x'�bt��Ɨ�/̲������T��Cy$�aVp�N�,��ՠW�(Y�"�zC�@a�����I�[8PÓ����>�*V+�Gχo�݁)U�P��1�J�����zk&j�(.h�V\��2��+!��>��m�*�O����rh3K�7�����M��.������d�8�/�p��[��s�%O�obIZE������z�j	�r)#�P{<J��)=
�E��q/��)�������m
&����6����n�H����ڬ����ln���-�&��W����>{t��p ��e�l�n��HÇ%�e����`��׺�z�^�`��˼	5[�����I�<5&$N�+��һ���ce�O!�Hu4�CVσ���,%��;�Ҵ(�O�۫bJ��T{l�E
6L����d��U�V�@i;gGeE�
���j�˼$��U����6q.t��ZL��7�u�V*f��W����Ȯ';&Up��c�"�)@�(E���<���n�@�l|��C�=�h ��Y�Xj)�[�'-گ�A���F�������ڄ�}D8���dN���ٓփ�}��\e�����2���~� �$}2��'����޾�ƻU_�%f"ww�;u��"2ѫ6L�3	���k~�%�r�s���� ��� �t���ϼ���4V�])��ߏ�]����`{�U�[A�z��w>��K-n�.p;��)])�!��)�L �@��B��s;�BΥ@�r�\�3��1:�T,���<���%ڑ�A:�ƚ"���ճ�B^ͺ�Bk��8�z��w�#��pX����Z��c�b�	�w���l9G��(E�Y���e�,��k~�ql.:�F}�
d� ��|&]Bi���3��r��%[��h���,�{��I���ß@c�TA~�R$��P4F��F�P!Y�i�����%���<�������^6
�ylO���xE��VV��P�� �{ե`����.�#DY���1!l��2�d,�<�T���d���fD�4���?�"}A5��v�GUt���?��D貛�n`�U�1�,Qzۢ��$A�*�]�U
]��C�R����y.���(�ud�K���(<������ɸyyu�>��=�(�#��B�'���ɝ5��H��Y����� ٝf�����|P����'�c_��u�mo](ۀ��YLV�)_:s=��8��C���JӸ�9v��@^^�%�:A�Z�9����a�l��{"�Gp�5вw�>*���ySӳ�|�t���t��89��<E�v�����KK)tx�#A�:��������vy����%,�B�i��AR��UL>ۗ�H��%K�]˭�gy;�؂��o#*�ƽQ�2j-'yd�3�(�3�W�XV����9(�wV?�(�M#�P���;�Q�����Ju�t��N.q���G�/����)��Z��J�2�0]Jn&�.f���w�0@�}Q{���Jj�����ھ��������Vb��`ы(�3�X�p�*��:�<�=U5ʛ�Z��OՎoOҞD�#��PM2�#	������$d}�/�8.:�'�ܬo�>F� Ȇ�8�0�A�ڽo���γT{l��+�r�@�Է���{��$�W96�\X0ߤ�c�_)��Vhkqf1�����#-����5w)������|b�7u�ӃP���j�TBBS��'��H�o�z��H%Q*9�uN#|�qKGR�|�I��vc'�#oF���q,n��dkm��H��ꨆ(�J]�^ ���Bg��-8|	b%,�e,:?�����O�kW#Y�f�8	g;��/!��
)���J�q�SP���~`%Km!�h�"<�>�L�z�dDd:�c���z����r=��:4F"�	�%t���C�=Ac�b+���A�PE��E`1r)g�״�D�X���)U,��x����y����TK���>H��C8�X�:녇����$������E�&�A�oX���O;��Q:�\*�k���TԷ�.���W.�c�u�~ه�fr�H����NߜY[
�Y$,�p~+�a�W��anC��y�E �U����m)d����T`���џ���V���y)c����t]&�tO�T[��r؃_�~�#0�T��8s��/I��;Y����@x ���7[�,���d�Pu����O(����h�&��Ն/��*���@
p,tZ �[k�n4���J���eL!+Q?5.��YÌ�+�\z�eSQ`-v�h��K�K�D�֋�J{!1a,Jh�҂/a@��a1G^���?��5�B8��{1��X�	��s����}"�4^}�/H?]�]�v,���;���u��,7�Ȇ�t��7Zw���.��=����G4̓�o�h���9���!�>�XS>s�dӤ7jy���������36������",/�݅ϟM��3(��V��2�k��[ ȷ��)�S���D6l�}�"�Yhwڻ*��GP�DiB�"��x�)\�e]H#>�-Hl?O;���q���gqh�����t���y
S���D��4M@��{����]7Ð�*�b<��j5Ҷ�#8YJ�������>�E�Wk�[@��jJ��CF7TH�w)��3�GB��"���������9�-�/Lq3|xG�fN0�A���K4�Q�}4�0�;&!_~Qͨ��E����|��p����{�=G���?5��8/�����F���s	B$����5��xUC���_�/�va�Wq����|+Jݳ�K^�;�B�6\z����\Q���u�{s�)���ť�g�n2�wM��u�'Ku�OWnK��W�����[T�Hk4���^b����E�Y2�.Zߍ����+�tꈊ[j�ǵ.���e��8�����^�|�ti�l`�ש��`�x�� �[�J̫�'����Ck��ih/���;�ړ+5P������M"y�0�ߊ�<x��e����A$�`��T��!�Kl� �%P�����*b��˞D�~�ol�#m�@��C�d��g��%-w`��i=���#I�d��P��Ǐ�@q�/�n~@>c]�'eZ�O>����� ��\����f{��^c��76�a�<H;��he���uqx���A�$S�4��8���N�ć(�I�0����W�<����S���%N��d���oMT�_��e@�}�F=h��?����F?h�PR��NX��T,�߃@�|��bي��gT�߬/��<<����:�v�Y�VX�s^h�.��́���v�c^��_��I�����h�U3
���&�t`�!���3�k��1��g	��p�����	�ź�i�T^M��6!��	IW�N����Q-�B���r	������B�@q�@��Ml_-��_��D��,���4-�z�]��|�>��\�px햾���kM@��+�٥�:<?��h�O,�+����Rc��ݑ:O�M��Ū����U�K��{Q��^�űxx� �	�V<�(��(�����Q�t�X�}9�%������rA�%� Pºg�$q #��IF"�o��t�T��)@觶�%qRv�d维��$������&[����X�<*��מ��zPˏ^QT�����P�QC�S�'[T\�..|���R�IHV��_lI���!�W]ĥ���OK���^�D$\� ؐK���	�|)�"��[��0�����>�
�\"�	�ZN���+���}E^���
�+��Q�fC��xV�f)�I)lsm�G0�
���:�)V�.y��Co�8�1廜<l�h�^E���^�j�L���i��~?�r�z<zß���%��:��6���F�,L���T���)�b������\�*	R_zWQ��~���2m�@����HH,[9�L=���/��A��]0�wA?��y݁hx���x�(f�3ׂ��U�'�Բw��-p����Åd�-����-�� �P���X`m��l��D�}���  ���3YEvPü8��V�|M��W�?�������G�*y��+��ǅ���?�v^�=�j���Yگ�d'gi�K�,Q&�1 |�������C��;��b�})^�cB��|�ō�Z[�6�o,��������b���l"�؋�E���b�)���rH`(�MV�{�a2�]OA)]���P��Zs|A��~뮼 t2���\���ŤB��~������v��A/�QN��RY.�u����v�#ʊ�@�����18{4Y���K��T�zC1�Śk	��� �߀W�(��IދF���`.*��UA١�jW��#��3<d=�,yS#u}�2ay��|)�(֚Jrp�W��j5J1$W�*뉟ߥ]���y�T����,�j�i`����G-�@镳񒇎�O��$^��U���}�k�֦.(z�%��zȽz+N��ޚ�*�g�k�)\K�'��M�I9�+
�Tj�0�uD=[	�Z�&�$t<��Y��S^y@�������U���|d�)�ja��(js�8Vc5�C�h�HEޮ�! 7�{i�h���.Z>��HC�W>���Nc�89Z�3��7YH���s�X}v*���t��#R����Δr��0����Ϝ�]@� �x����]�};��q#�U�9j���ױ^��
3$�[�ܒ��@ON�y _bTF��ʽ���>ʹ� >��v����XZ�2�T��+��nea�zT~�	�#�R�܊���:�J0��Lw7.�DfUi�����ek���Q}F)>��e8�X�"��dX���<4O��H�-��Z�J�Jݏ���ɵa(X2^�S����u�X�����"I4$�|��E��3H�*ܓ6���"N;��<��X�xU����V@��ѱd�\J�j0\n)�@�Gh��i���ԩl̟�V���`~�b�DUw�z �h�����ÿ ������p��1Lqڂ)�CA�k?J�pڿ�ga
T�[���M!HR�h��[�P��$��k�T��x���JQkS����1�]X�$n,'��Q-�������y�TN2i����]��YP�[�bT��&�9�b�B=w���玚�G�Qr:W�+@���W$��ŬZsK�P�H�Cv1*R�Q%���\�2n�0wK(E���!@�I�j'�{(�z����#���5�N_Tp^Q����R�z�
@������G� [����ɹb�OZce���/�����	U�x;7�CzG��)�j0�R�S䞮G���^��-�{��!((��L�K��9V�Q����Xh�m�P�YX{<��JB��O.�IFZ��u�\�����ڦ�@��3��)�0���@g��3�����s�*�BNS�Xܐ�I^�!�z�he�$t�7�z��T���ڕ���h�:�a�_	����
����V�h�^�ȃiq�ml=�����������",�r�M�:>˂p�*U�r,�W�����w��0���@�������R�³S��8�B�!����z�U�����Q�b.<8��SX	^�S�=2���lS��j�2g�ŜRr�e;/�^J�YW�q}���5���^�ޜ��FI�s;��:�A�TV(l>�j�U��Eϒ����
��JDr��hWx.�L�εZ�Hzw[+��J�_����{�҃<AsI9�n�ߪ��|}L��v�Wj-N5�n���;c�I�)Oh���\������H��U���{�L i��|Ws��D1��e�����ҿ��_&�e�}��I~�_�T��|ʊ�V~��^�����$Zx%��n�z�J���ͽ�h<0�d��@�bМ�+�s����wу%��Ef}0�aV���FqE�JH��r�o��u�}�~=��	XL��dy�^g ��l�ob�۬������\Fh$���T���QǴ���Bt�E^r��S��i��W������y+οyVˮ',���v.���V� ��T�x��\�hg6��\~�u�j����Ti�+�������G3.؆�D�ݨğ����͐y=�������un-C�-�����t�zΊ��(92��RhZp���)�JH58\�@�ӹ׽�(����(��$r���h�n!&��m���n�T�m�շ
0�"����b-	�4]6��p(�9y�%����d�}�I�R��LѮ<}{�.FE��f��D�2�N ���6.��f|O"ÿZsUs�����$���ݷr!�\��H��y�C���+5ğ�Ѝ��Z�]c��5<���S�I!)���;���K{;ڿ������%��Dz��"_k�C���n?��%��u{�&qB- ����ۖ�aC0Q?� ��N�����[���NeڇI�qˮ8�[��]:Dt~"���PB5C\@�A�)sM�-2��n���8��qV��d�	?�']�������w5| �z)z�d�o�tc�Ok�V�����!
MBx3}q*�XB�]����������ޤ_��[�a�a�����>ٽ��*P%('UD���� �.>`��
|���h��b68�H%A����Gvr�q
��V� !��Zt�~���v��g�|��hQ!�� ��x�!3���̓F2��k������s�Y�f��e"���'��H����i4g5y��^`�������u�3' �����5�&=��&j�~O�kB�`���kA������x�"�M�[���	Q�h�c���^����xQQ�VO��_[	mg�4f��Q�{6���)��+$�O�������cݼS�W�\��5�Z9Y㥝�xd>�����X��m�nT�1�s�l ��d@|���>�q�e��Z'OR��$b�;��Up�4�/^Z��\O�&�|R�+Y����Z�!�|K�T�j���W6�i�9�s����Z�;A� �1�6�!	�~9KU�����|��S�`�8����a2�HBt9��� �2D��,ׇ5dYB)~�z�H�����ނ�WkT|L�G#����}��G�6m�Ⱥ��ȝ�[���+	N��/Ҋ��������5֋>�w;>~�/��vq�F��q-�������7±ص�Zۗ��f!H����Yy'�s�Yny���S�ez <��F
A˰��d��-�Z��Z�"k��k�e�|�Č��-``�*�r�+�뎏!��Zj�o%�!}�����^Q�E*����i�Y�5 A��$��BHG�K�?�U��P7�Q��~�m`e��!Ux��V����{�u��p�)�䮇����}[��c����vg��֚%�jZ��շtnb�0�:ĠW��6�I�3t;��4��B%��ԛ��t�U;��ɹ���-�+4������>�F?��}����5}��Q^e)�[>��_��YR%,�`;C�*�~�\*����9�O�$����+�������i/�؞��r!�ɓbߓ)d�9ci 	��|
gvi�#��T�	^Mo�F ���-oA�(:�!W�FX��PG�~��ZmFI����ϴ��sm�4�֡'��z� �R4,i��	�w��F���?9�\��F=٘�9Z?��㬉�� ��M5JNB���?���
���m����~�"*F�E��S�iB���"�u�[ĸ�*��Q�"��|�)"BU�ECp)R�BŸf��"�����{^�μɼ�w��{�9�{��G�>�a_�^��>ʯJ�}5=�jZa*����i�{=��!��g�I ��a�l��pt�'m!��U�<lg"d���3��ݚ�7ص2��2kpr���<B[�E�����R�Ǔ��A.��$�ar�r�%��Kk���v����*�`�Jy��mIkK>��d�b!0��zO�]&�ԕs0��0m�UU>�CO1&o����,�T@�\×�=
;u�kQ�'+щ}P��A��L�:��y,`�>Aw���e�t�|�s+g�ɨ~�_��)w�(�P+B�J��/���:��_��tZˢKY��1Y�Y�ݾ�o�d�u -o�f���r`����nWv-F��a��;��[Q� [�L�;�G��^�J��;
�6%���&;P�]���l�������Ҏ�kF�2���9*�n�^[�Z�O��Q~����0�<����JC�% �3hxn�&� �cm;�
��1V`�\U�Ci�ʺ���j�M�w�߀˰��P��FQa D�a
�bN��{9��-��ت�������������\y<�d2w_{�_lGi%�����f���.v�j��b�ݸ ,N���R&������~��9����?�=p�v�{:H9;�[:Я�h��a�^���x�:~��Ý�y��֬R�r&�zف�[ٴ�?�|���{X�7�_6Su7e]�
އ}�K�
����Ë�%U^D;��tb�ņ�������tT����6���p�d����НN'�U��6��Jw'Yw{|�Yeq:ci"�;ͤ�k��>vd7�m.���;}�4����R
o��4��鶸����������s����`�*��J�YU۔�����Ï�ɝ��\�w��GnIy�+����oL�����e屟Ƶn�h�3.U{�	� 	�f�Q�?����p-��N\1#��;�](4B�A	��H˧m��wC�w���Jl���>|��5�nh6ݕX{�aMm�[Տ�1/��~j�2h������b�|�5ݱ�gA�F~̳�Hs��"W����0/g�����W�L�஑=p6N�G|6�y8�~�^G�(����ap ���ԫ�F����G�uh��l g��B��:��H�|��R�~~ȐYo�t��������reN��ʬp�6�"��� VI�R^��h��^VI���_;"��)��kG�y`��Y�G:��K3M�n|ن2U��ZO�>�@�B��ņqm8�ƈ*,�ƘŌ}�-�^>_ƭE
M3��C��Q�+fR&��T؉r�iV���a��·+�|�����Q��sQ�3�T�\�7�||��^�6P�23��F���7��h�`�������<G7i�V:UyT{@Z�ɥ�Q�T�)7�BD�b�n�ޮ��X���
v��c ��n�`�>ǗB[oa�;a���/��zþyՃ��N.��_ѝ^����=���	�J/�FX���:����˟Ӄ�o2�~�i�-�����
o�e�e�*��E���"�w����	!�1��a���;��`c��=�R�o,��徼\�*8�� `K���W�6�Yɥ�]�F�mw�g��?���(���
v�ng�(�C	#ډٖ���i��rLu�܉�:7/�a� �eY���~K���@��N唐Xů���HV���K�u�f�p�>�3,�b=�uB��Xu������
�9���B��"1V�5��-�.AO	[��_C����E�b��ڄ�0Ϻ��:+��f��jo�o����3�+�̻��W'H�ze�Y�z�������NX=i/?�򷚤1�
bM����Q�8G�(�m����wٶ��	�� ������YE�E���Ky��8sT:�:d�u������Ws'oW�)���߷���ӌ��E�ɾ����tq@7�t(V���n�  ���ǎϑ��yO�}a��J)N��<�1r�M�`��I��d��vsd� �H��}�3���#o�~��!�5=kr���|�4�b_ɥ=�?]Y�[�h���m�aJ4M@�7C��Y��{�4���=* c��"��հk����L���V �z�D�����d�9�?���f2��:�Tp�x`Jrj
�F�O7���S+0�Gﵖ䣃..4bJ6oc�"8@�W��ۤ�
6�W����_	�L��c�\SQ�3��w���]/n�ۡ�5u"����]`a�O
�j���9��?$9\a)��'H+6/��5��*�l!Rn��h� 2������I�/��
��^�*4��}�	�o�9�K	����]�(������y'�|��I��L����'��of�o	;=�?�]m�/qԁj�UOK�K���h��� �(�Q�N�hzDp���p�U����0�9��7zf���~jlx��N��1������pIݩ�i�&��+Ŀ�x�͓8'���-!ՠ&8��Q�S^��|�P~9CP>��Ey�_�xS�MAe��K�wp��t�	���M����ǳu�߀�����)zPҾ�5K���I�:��0薈�����?�S&�(ahk�B�4��a+�6/�0Ql��J� ��h�A�s�e��T�
S�%,L���~��nx���"�
I�3+�i��i���ֹ�!~�?�l�^�q�����ԋ�ӂ[����A����ͪw]��=�B�dѿ�7���>��BD����6���b=�z3��w^�;J�=(_J�㣎�W���y��,KF�r�����d��BI��i��S�{�y�d��Uz<}8k\�����!�`fȇ�5L�
e>�qH����k���=�|ӭ/�j�X����D�s���X[
&'�1�_� "��G�W�;�lTO�~�<Y��r ؟.����Zi:� 4&��J����"*��z�{9��N���.甐�����D�i ��+��˘�`_c�+�Y�zI6������=?�:�I,� �V�_�E��������:�O�s�G�%u������Ut����ȧmê���g�î��99T�
�I�`^�������@��a
������+c����[���'�F9�#��r�W8��Ю�]ݽ�,���KǴ-�a��^o�Z�Z������R�IP�PO�����b��B�<�Ȗ:*M�}��c��Š=i��{�ɕ'^����I��\`�r&����~Az��Im����l^��㒴�5n9a�]i^���ݥ�cJ%����ԝ���m�m�r-I��,�4��e��H�`gV��@�J�b��]��r�$y�y�w�a;P�Pka{u��^�8�1��0�`��8�y�� �h��~N��J~ �%�,����cD	��[�I�]+�m{hrK����&k����:�J��vZ��a�_�5��L�L`[�w&�'�ҹ�v�,���9c��Q��k7�Lw����nE�`������D�v ���upc	��\l�2
u��Yl$u�7�,�;Y�3`� ��K�����]����z)^OZ���]�;���dW)v�L�g�3o�0�| K��̾�?�g@s���A�.p�n^�{��sZ:�MD����C=�ۏ|���F~�Y"i��T8��c�:�.�a.�ڳ��\��~�Vg�a�9��b�k�	����yĊ�mi�����Ka�:s�d�X�g5*���:%f�2��b��2��qvנ����b��Ls]b���'�1�6��Z-'���D�Ӯ7���g�w~K/.�JCj�5d��7�� �K��(SC�m��,3�	r5�ȹ|�FOŘ�7�<9@�/�g0����|$-�� � ��/϶1�� ��6,�P��г�&��eM=�\I�~�/�Ԯ���W�5�gv+�1�~����<0b�w�#��Z����'m�����ķZG+��.1'���'>���C�^��<ꗰ�Ft%"���qq~1����+�~�!��M���e��&�iG0��R�#�[C.9���;%�^���C�c�']���+�e�5�c<D�7��2:�����:�,��״�������:o�G�1��γ�ʔ��2~]��ق��"���^� au�AΟ����l��jS/7�Bī��˘��aS�a��A/?�l����3 �5��-|C�Cr,$]�!��F����� �3)�]���4}�a�t�t�eB�����VU-� �~��5�0"%zJu�OI�e�T����Y����=)�VKtAJ���!%��<�r��-X��6g�x��0x����ﺉBy3$��2�%��M��J�m
B	�C#g���\�`MW�A3.v���,RE5B�0s�@H��0���K��cT��F�}��� �լ&S9%`��̦^AP\ʬ�Qt��g{8�Y�{��X}��P*�	��{Ȯ��l�'�nC���\�7vsIǍÕ*Q�.�ձҐ5����,�����OSGiO�#	n��i2�1G�l�r&�/W���I=UZ8f�F��\_��R�G����V�P�K��&���TYB5��i��^��������/No͑T�Ũ���5��r:�Qz�{�U)Rk|�}�r����&�:�i��U_�3�߃���d֮�f'��9�?�-�*�����^��E��V"C�G��W��C�$�5�h�83�Gi��@���|��ϔ\�}�v��h�'\-%gn��+
���I
?�.<M�^�JK��Od��� ������ ���tV�ű�B̊�}�)� =O\꣜ALه��z].I�=�+���8
�P�.iDxU����  �K���GG�π�E�6@����O�k��Iuͼ2_����(ٸr.���Aʧe�yOY��iB�Z��IL�ܟ���7ј�8��Z|������A��4��G���̡�0�c�����I�ˏ��{�˕���j C�y;~M��� ��>�~�&|��_�x�L��7R�Jʉ�5A�~$�r���W��Q�q�b��~zl��[H��Ov`��|�֕/�;r�R�p�o;A$+�j�7�m��<�|V�^#ǡ�Ki���p��V[���3�_�N�2�\�_�+�t���Mv���X�ཞ�r�� _���"'��Cru��Qއ}k�0[J��9I�p�x�#-�����%�\"o����G�� �3Ǣ���{�m�oٺX�X���%�O=��#@����K�d�5H��h�����Z���".ĊH{(���������!p;��R�Ό�P5��)�f�r��wy:��.�y�ᮃmv8Br��GsW��e)C�:��R8�]�n��S�ڊ��y��zc�����T�܉�.�"��x�k^�ʊ�5?�CV�yG:z���c�,ԫ��-�k��0#E�$U�ܲ��hT�-��{$�|�����w*��n�X�؟�K�O�<�s=����&��?�Ӗ�:�?��y����K�2�W������sL�)�,�D�^�_y0�ۓ�۸���h�t$eZE,�+Â����_h����&���O�)qEr�-b��̔�ZV���k�/�{�i0��ǹ�s�'����E7;`��:N��2s[��U���z�J���_L��ك��-�� �l{To��
>�@�Lv|u�o��p�l��ndb��~X�ܝ���ҟ���{�;Ճq����᧴➦�Kp*a�N�nU��hx����$����җ:ˡ�4�T�89טl������b+}d!��J��m�;.�:Eh���T��˜}�V�v-4|���)_�����5�s\��չs�� �#�(K�8�1����m�A�+������>S��� �$���t�j��ؤ����|��8����;��,���z�W�j˨K�ϣi���*�(�;06��B;�U.�w0/W"W������R+B�+����[ �����x����T����,�ã�&�����0���WP�I�\��}n��ޡa�@�"RC� �U�0�|7L�Q1E���8%"~{/���
��:��2LDfC�#%�=�!�I���C0MU_��=�	W�a �V4��]}oE��J^�נ��`�NS��A�i�	�aW|��ŹA�2�G2�CN���V&S�?K�ə��8'�i�TA�G�(���P��gX��a�dX�}���~^�/1������e���2{Pze���O	��hC��r��K'����>�͌��oz���8d/�e4V8��F���v@�}L�X�T�ͦ����
�^S=r$��_r2@	�������˝a�cM�>T�Or�-&��4��~i����D�B���Q���QM(����r�\*�&�u�y({���Y���(��ޞ�\Q���y�q:�5�t���D?2߶��>b {�$fӉ�t�q�J�����=D���`����J��)���.O������IIW�;ڤ}����k��o�r�ΝX��2����i��	�t��S}��Ď��¡��z8&J��[�<ݨ���(��{�'�Mr%���0.5�'�Pޛ~A7=����� R(�&�|J��C}\������"����Ky#���3����~�E��-���Ǯ�>զa�7�:^r�56b{���{R�����
r+�5����<��0iuq���nU����N���S���W0�y�zS�}6�%���:�/���r�'��x�
,DP$|�59�,��)�=*��CHo��Ĺ�}+��1�(M�ًe��H<�
�QL��H�R�,�<��j:Ƣ����R�1��鍞��B�1�O�_���t��*w�3dy�9��Mӵ�5��z9đ�v9�� jy6�
B�,v�%������C)I��IB���"N��y�t��0�l��!�j����<��gP�~����(�:���H�X)��i� P�RF|�b�l����Z.>YY��243"��>������E	~a���������}߁�}����{�9�{���s���\s�դ�#G`h��K�ڿ�2���{�H�)5�j��9�eh�2��5����,Hod�i���e��o���l�cz/�	'No��ݓ$�fSo���Ia�>1I7|�RK<���1҈�����Q<�����B��$�}��XoB#���ЇFl�[��@h��K3to���?-}'�w4�b[���A�'�7�	'_�8 ��S��_F3̬�Bp��M�P�޳;�Ыs��μ���*c�o9�k��Cp�ԛ�~�Ʋ*Q���:GAA�Ł?�m1 �*6C�(�'<kd����'^�м���A	��It=����k}K�.�?#у�w?�q�+a+ڽ�bv�ț�^�ӷ'	9�O:Z�t�|%���8��Jt����q�;_��V}t�K��zC���<!��P������N��Fܕ�#T�����d��oЪȟ��+�ǥ?�;1��5^��An�_)ދu��-��9͒��ظyx�j�}�K�Nx�,k|�̸��O��x<�1�*�h^~YQPt�8�~?�z	�W��nү����0�܅D�4�}��K���>э]g��y��?�]C��u�q'�X��K-��*K�<���)<o�Y!�Sȹ�`�7�m�h�t���r���:���|l����6�~[7�5����P��}�L�5YM�'-�c�d~����X�Ht:��V���G�#�}�4���Y��MD�&g��j�:-{G�N�a����3+��a����s��a �*�>V�ET7:�����N����l�w8��������x�	j��B.Ҹ�����)��^1��F!og�}S�X���_��ƫ.|��x��3��BSx�;]?}޲ԧ� �lώ�O��̦�)�M�����~�U��G��WZ��g��hZ�W��ii���u$^杯vʪM1��ol��6K^�]�J�K�ݳ����ݨn�ŵ���ܹ�K._��\
�Oy�r#t �仂��'�v�s~�/��?g�Jr�E��$"@���tƻ$��Jr�{������ � ,��0 � I��6Fc"�uo�u���&�A��O�f�`�X8*�z��Z�m׵�0�$��=f�n���tfq�����$KG�3uk�(�����kVEs��h?�@C�/�p�ӅٱȦ$��)ޣ�W��B��E��S9�H�\�c8V� #G��������4=�`](7���<<��4
ct=�z�N��Y��ʱ�ͷr���#l+сAa�ހ��y�e��+�U�N��D]+f���S�mn��(��Y������q�<c��0�"j�)��y0�T6�����h���A�d�S��-�MFQԋ���r�O\E�"�g#��H�"�������;�f���S���*3��l8�qr�g���3r��iϢ���R؜؁����]� �,p2Dj,|��zR$�l���!��$�e�nFC�L1tc�X$�����Is���`�(r5?�;6�QR��.��K0j4�[!��	�!�Я'+ѩ�*��]�H��'밋>0�O1�U��Z.���A܋��uC�>&�3Ɉ�V_*
cz���d��<�ȍ���:u#��A����Y2b$~��5I<�~0�G�eغ�P=f��������cYV#�r�+�������4�>�*��4�f��n`8B=��9X���]Z	��H����� >�}�e3�.)���6��hKĳ͗�k|[5�M��j�
,$9D�¶%$���j��$��|=���l��.n6�Q������|����m��p��\��3���B�֞���`�y�C�����JǨ�+��!%�}�|��L�j�ro~[����c��M����Z��	�Q�7m���� �����%i�P�� ,6S��6���F�:�,}��ˢl�	r�����7��4��z<����q�c�-R�]0���������OP,Cy;�_��n��[����(�7����m�vk^��h�H�!L��,V�\�M��"c6s�T�W=��)�S�dU�dFҳ�+qD���;*5�1A"� �Z�t�W֡�N}|�+i��I�4Uέ�;��pڀ�����h{������ԃ��-qƅf'dx&��2	<	����-��`R�`(Qxy�Ю��x�z������bi�7�~��aqॢ>"��+4 �&1(<���R3_�o�����p���ó�u�-1J�r�q��"��-,;�+������Uh��j��_�����NBBc.3ڟ.=�R;UŐƮd�xX'a�
�o���ڿ	12Ҿ��qb�ҍ_B�;A�`@�e��1���҈�c�хh����lЁo�[ �{Tn�NGs�kYyȂ�f�C��)�I��S/����Q2T�ۈ�|���n7��n��Po�>E�֟�?-gػ-!�q'5�6Bio���b�� `�R6�M�,0����u���bFs#�7>��%�g@ˇ~Axz��Pi����3����J�Ôw�۟���Ѓ]A��'�⏊l�3���~NB������]d��,Qv�>�"҉g�K��Ŏ�b�]}�2�ƌ{U�tF�9Q�ĵԤ����aU���H��z�᝗AnWikI=���CV����p;�wY�TVQX"�b8߫ω��h\g����s�f�ـ#������[ ����8_Dw1+g�F@Ҕŕ�p*4�Uʃ�~��ِi�)
QO���2��!ml�^/�h�!���46����L�E���ȮKfH>��j�Q[쓲f͒�n�m,0H����&K�`H-��������a��z\).���ϣ$��c}�	�EZt(�3�G��09���}Z�b�:?Gdh�����0R��/�Ro�|7�l0��Z�ٸ1�Y�J����h����0�j;�Ӣv��=��J�|x�E7;c�r�	R�ۃ��0$�jM�O��e��đo#ܛ�b��'�N�� p�K���ڻ�-ҍ��ƙJ�y�:�"l���ce��tsl�h�FJ�� �l@vbh�F����O6�',�=@I�3�~�OX]�Lk�=�gt���1{g�l[�-�J�Ml'����w}fY�ó���v�o6|Mo+]	�ߤ�����^)���?��e������_���� �QaB%<�|L� ���'��CR�9��%G�<�}�h�Ty�`}��^�I)�������;�_�)�e5������P���ȣasx��O�ؠ8���nF�'���p�x��*�l[Z���+�?��Si�321����΍�Za+dd�gc�׌~,��^���F�,��'@7�gU�?$����_��e��ܦz��~����N��#��M�\��2���
�w�Ŝ�)�(�9/Y��U9�����F�{XȽi_gd}�
����!���k��G Y��ی���E|���L���uغ<�j��e�eQߗY�"؄�P3�,M$�8���Iam���
������ż�����{(iU�����q�Za8s�0���#�a�Y^`������h�����o�x�o�ɜk�G�l�K��ù��k�,F��#�08�3��DɁ4|`�����>�J���7~(�����B���"�D-���a�cIzYd�����ŵ]��BO�Lr��k�h}mP_�k��yã��ҽpޘ"q�q7E*���_Yq��;��0~=?�������P����������01~���i�\A�B��7H�9�k�ǳ)�lPB������K�1���Bh���@���Gg�,�w����^��Z�����ʍ��¬���s{��n��m8|�*�������6Bz"�S��aw4g¾���.�ϙ(��1����Gy�Ӆa���+��<��<Wayem�	��[[V�k��(�ط@���������r�����Ѽ7Y#1���v/�u7|/��ď������&�K��s�.c����elg`�ro�/�.c�j����G�p�Z.T� &����=�O3v��`ay�~���]�\f��;��ˮ�p���q��.�+>��y����)sZM��Z�����I�K�z�|��,��oeXW|8�J�`�
~�@�7���p��)>�0�����&���T>�[�'��]Xͣ��L�}�޴�[MQ�N�w����1Y�<�4���o�ϲv�>��ν��#�sB��7����/��S�N������N_D�1��)��U,p���]n��K��7Yc1O��ھz/E����j3O]�#���0}p��o�>^O"�)v������ey^�O�:d�)�������5}��Y�������O��N9��}P����l�@���2��T|��-��^��3聬���j��wA�rt�˱�}�V��-s9"�'*� ��^ix8v��\��H��Ӿ�r�h�I>t9^�1�����8�d�GY{��W-�%&����>�ll��k�p��6Z�u�����q�5������d������Nͤ�q�I�gg�a/�4�uo,�=i����'sMO�5��'�*cǏ4)�W����F�߭����qE��C��w`�SѾ7�F~���v�)zp6�qӳ��I>�$S��&�M�tg� \�'g�"ݜ�������CJrI�N
���<�����S`7�]Y;y+k�d�\�nTݞ���,s6v[���&;̩0A{<N܉�J��ӫ��U>Ƅ=�'�w��I_�YwN�Hkw	�	���ޞ��R�����#��ld��	�^E���(X��_@{��tY����; ���"l3�>�-�|?�Msf_�z5�Q)�&�&�w����Ջ�X�Z@'�i��b�,\;��F���UF�IZ+GZc,�碱#[@?�2��tR�#���^X@_��PFY7�=�ڐ�����p�{���-�tQ��~�,�]�K�Ѭ��~���¯KE���V$v��>j���`�R:�s�ېN��֪��vhW!�v�����hÖ��Va-����4pu��d�n�hU�RX���L��I�ł�_6�<F���t�e����*��IfI�Z^��X�Ʀ>F�TڱHu4�
-ʬ�+��`�g;� L��d��$f���A�a���W��Q�#�`��Ѣ>&^�Cby%�'���r��Z�+�(�V����Q`�]�ˍ}�uw5_5 �`KlU�<.>Wz��Ȥ�`/TF��i6����iZ:�#�����d)-|��:�(Y�4�H<����� ����w�	2���g�| N_��#\�=���g��%�@ɥ�w�a}+ot�?��>+���)�C��݈K�D���0l1OcX'f	2c (�p�������� ��2v����7D@]F��0;��*�B��}k#��t/r�Fɲ���_p
�e�X������x�#~�t��ä/��ĺ��?��OD��f�����G�G�O�aY��7���Tl�P�q~Z�q���)M���c����6�䛳c��{�E7��	ߕ�˘��|Ao  �^��̤�e��JA�ˮ'gݕv�:lZ���,J��I%�?ت��4lt'�D��SG���B��[���(0n|���Q��A��[&�PQ�1Cŗ��D<��5�{߀�x�O��t۬�<P>ؔw�#V�t�a`m��eO«����ֶ�K�x����;w��~����K��Ip�n�~��S�X�Z�bqZ��W�}���`� {ͺ��7l��|d��H{9�zq߲	�k��j��)Gs��}9��5Vp�/Gl�rtG�����?�Rץ]�Ƽ˻X��j��k�0�A��
�'U������f��/�����Eňtg��)#m8-$�k_f}���
���F�U�ւ�Q��:AzK�kM&U��
����2wP*���a>G{�Z����L&��_MOw1��v�$E�j�x�f�]jF���Qvk��mXn� 2��Ht�Yc��Z��'�Kw��*�>U8�"�_�Qu��I͝G�ק�N�����c����]��te�����Ƃ��;����z��^/
���w>?ÔswO�o!��2��4����`����	
P���v������6f�Ji;�h�m�2����{<\��~�	{�5e$�����>��M��nQ�.�1�}���W'���Ʋ���U�Z#iVy'u��D`�ജ$E�Q�L���ST�l/��kݕ��a���"#ۆ~���qD᜴d0~�ʤZ/ޫ�"��ΐs�M��t�³j������4�O��#��)�iϵ6�䘌rn�c���Y;�p�e�<�=.k��G��
��g#Fko�vk,'w����h��'б��ru��L�wa���֑Ku7|]�]�k�������t���m��v��G.C���L���pn懱KSl����� >>�8��O|i񩲟X�nc�O�se?q����'�+e?�?�s�{h�Ѧ��p�6�j������.�vF���� .gd�1�>kJ�N���^��\�M�	u��B}28T�k�kه2T���� v����J1�+#�F�KRT��ji�ߛ���H�����,�2&f .�d 9|1(HrNP�2��R� 5�o��5�>��j�_���}S� 1�{g�-|؉�.�|\J�S0�b[QP��pwI?��̌�ִ��R ��)d�U�`RPxb�LVo����*�Th��yM��ؖ}8<�vD֍�F�@�g2�׍@AnWd �!�J
u��Z{��z�����o1���D�)@,@��	���)G�ڳ�g�2kzL�N������?V���|V�-0�4rk
�z�8��/C�;S���L%
 Od*Q �)�[���Mi�]���OQ^98E��M�!���y�n�Q.t=1(p1%(��@A�s2��X�F���Ge #R��j�([A(��jL�ߑ�G�/���0�)���� ������K�����(?Ț6�V��/�?}/L���lK�U`��f/T�$ㅡ�~y��[ �k`���ؗ��vX���ά:b�~�M%٫B�����oļ��I�Eh�����)Iޏ?��GIvU��$���j`/XR3�R�����m�oN���Q�ӄjZ�$'����Q'W�(� �'Ir\>U��:m�#IvTK҃��S�F�_���tr�M�8'@|£�������*�h���pj*��ڔ��X�D��K��zdvėJ
ax�(AFT�6�a�������Qf��AFeuL�a��Z�'��5�RSk�|>�y��{��������;�w��<�y��������&5�Zo����R���UV���5�H`�
ބGG$5߰
��/�x́R�?�t|R����p�+����±E��Dټ�K
�E�n�|�Ҿّp	�K��yI����+I97����ss�������J9g�%(LS5F��"�o�IM	��ε'��`D0�j'6& ��L(��:MjN�6 #���,�,��};FA.�ʫ�mx��c!�6;|��/�`���h�T��#��+�[=�Bﰏ-X��QЉ�泚�e�*�Ќb�HM�8�(��o����t�݉t�"��{pu&7S�g�u<k5	�(��}D��F�G��WI���Q�-!�`|)�H�w����{�I�Y�)k>�tk2H��c�ꧻj�O�T�褛|I%gf(�*a8Mw?)�A�,�%��ҁͥ��Ч��y^@E�e�ؖ;�*F�/���� %��d�M��������'�|��푦�xa3
�é7?'� �~+�*2w�Iǝ?;��Ģj􋢣O:����	��`,��4��<������IOK�������j:���x�tN
�h����X �Cl�rZ��I9-�[�rf���5�wI��n��q��o�O%��$��a�8��ٯ�����tr"���Vd(�Iyd�#�o���Aʐ�+�P�7	j%��R�,⯵¢�	̈́��`T�\��䬐&.�ECf��j{R��qqF�sS�=>��aM��36��6
)S�>.���v��'T�;r}Ȗ����33l9>'Iynr�g7�h��G�����Z���Ğ�+�ga��O.�eC�zƾګ&#��-�]s�V9b��w4�h2�f���,<���T�QT�#3�ԅr���r��jI�Y_i�y�g���;��T{�T�e�Z�W3�H.�S��e"PW�6)����������9?�
�9+5��g��eV��H<]-Yw��x�?q#k������<3a�
g<�(�t���}gP%����q��G�|��C��$	����	X2�[�+����q��޺*���Ǹk�:ƑIGyLR���3�\-�(��¿���	#�F�c9g�g����F&�ʣ��(��/Eqd��&̏��1��]�}��Z�Z~2�Ŏ"k�½F�s�h瘝�6dMR≯�/E{�	+��E1Q�V��}Q�5E���h�}\�
C`s�7݃:_���j����t{��W����.=9����G|Q��azB.5e&)*�Q�7,��6���N���s�I�?�K�_I��<��D��t5���{����L�,�q����z�;Iy4�իb�(#�P>Qd�$�4A&��?�5Y7�V���5)gR�ۥ����Ej�LH]�~҅v�ъ�K!:��n����`�mܪpߒ1�^sIȁ�P��n|�FzM�Fz+꠆� ai���9$+��������k�su����`�r�� z�~|Kh[ �;�nbn2�-�nj?�0j�1���^���0""�נ�ۡ�'9V FSC.������ѳ��ق�N_L��e�h�*����	o���(]`8�^'�~�bJ7���!?j��FҨ1\,~	��H�;`�;@�{�]T�d��s�Q��X���:���hrq���yJ��7���X���r�B t�CC�*B��/B7 ����PCWg��v�i�4�u`��B��`4��Y�B?)2W$U9]�s�\�]>�u���R�q�Xԧ�mQ��c3LA�Hi+)�y��;/y�31$u�4��'�ќ��ك 4�cDjmK�7��F�J����*aRļD?��P�@!0f~��(ߗ�2m����P�OC�eə��ZN	]��$��>��� ����;�,���a�PF�B�Ҧ�d՚]�A�Hg�]��E�Pе`�Z��[��b5�jk���#��Mj�Q���Q�*{#t R���b^3���wHJ4����tWҐ�s�;�����
##��<<�2��8��#��¹_\�Bۓ�$I�o�	N�?&�5vC���;Ra����F����H������`��F����퀈����_��T�Db۝�s�q��������(؉ʎn �������V�m��8��r����!����H�%H���'�Ru�؉i�[Ez����\�JԵ��L�&�y!z�GM�5�����B��i�X�D�<�U�v���v���l¾bg)%�B�j"Vn{yL���W(�&*
R�O(쁻�kX=���l�аE(l�`$�A16�aA�pH�ڐ�;`�)����e|����mz�Kv��4궷��y�)�e��E��ɥ��y	��axH�� �2�UMᐐ���@p
��A|�j
�&���B��O!��2
��1�j
ϗ�":���P)�m"�fz#�
7�R~~���#�B7�p|.H� ��ϳ:�����|2�#��?�,U��1�o��'"�N���T�zϬ��o�D奈
�����a�n������^��4N�?����O�n�w�ϰ	;�}��c�-�� F��>��*���5�פ��m�ƿ�@U�=�������;1���9�O�D�ȭ��2&V��G��7ľ�v�֚�I�/����ּ5i~D�X�%I��LsM��>�]� *ϻ5�?X�3����ݨ��3��~�]ʵ�\0�T�����Ok������/Z��P�{�{���$p�Yy=B����[��=�glu�i�W��\и>�ج�[�9�r�HA�'�z�r�0��(��	���ؗA� A�c��ba�u��d`>��Rɞ('e���a89�������*��20�E�ٳ�*%d_����ɾCP4!d7�����3fڅs�.�-����"�&�]�L�����O�>'��#�% �c*q~��b��Ǎ<�L���^!�M��1���]�M�)�+��c/���i�J�������)�N�p�E�9���[^ʽ����������6\�ϳ��[jP�?��R��sT��`��%E�OO5��wM�ݱ� #�=���ی�;;� �����`�+0���JG�f����2�Q�U�}��Q�����u����7XZ�'�dP�MPPOC�;��ދ:*Y2��"���x2�|�6�-��84b�~�6�`nv穌9�G�NN
����U�����K�sz�n,Bq)Ȼ�H
g�Ke�uJ8sb�wez1�
�l��
���>!gj@|�{>�bV�3'
���ș�3(ޖ�ţ�0��yr��I�|�(pQQ��A�(���3�
�yb�z��:��f��|�)���1������ׅ�:�,���v��b��M����L8F�̫BН�VaN��<*�~	���2�>�pz#�V�a�E����0�t$��!��p����y�^�KD92/ʳ2<y�JپS�(?���B������"hyŊE�����["�IEN� �+�]��7cbb���-E�)�rb���K�{A���Ӿ�(��������VgPȈi;>�ӛ����:λ���~-
�N���^�����X���ma2�n$����4�'����(�-v�)0y��p�~�d`WWdP�f("���Y7]ٺQ����a�v������7.��}�_��?-#���!y�>/�.��|*I���i��
L*�a�ˑ(����Q�d���HgNQ�v���&!�k�֜�؇�@G���37�� ��Z�*%��3�o�<���3��6wA|�ՈQU��R����\�B? �Zh(ޝA����,(�᯽�e��X���xX���Lo�*�ed�SX�r=�3s���a�$0��\#~��Ezr��R?S=�QP0w?�)1�2��M����w��9sL��30C�������4<C�}���I��KSB5���J�yBOx���OX��9������X/Ƈ�[�a��D]'�{Ƚ8aY`�:'�\l�);"�� Y�	�~�@y6x�"��`��ey䅿h��X�?�|�tɼ794>��b�8Sѻ�^O
[�r�mz��,�m�J�� ��i�ݛ�{��~�ŭ�%6#W�U��bLZ��ErquzaN�:-�,�ȺW�*̋�kL�����ϒ�ˠX*�:�G	
�ε?b�+=����1'-������	�Pf��X�E5�:Dv�
�yR^Q�	�)?���dMu�qU���L�H�2�x3l��� �O��R�	��E1��2Ho�n!��ir�l# ��IB�+���ѓi����� �#����)�[$�%6=	zî��.��.a�톷��r4�	�ً�ņp9�.(��W�9.��|�X�X���&Q�Dz�����`0��86y��i���Y��C<O}�a��q�Fu�V��[$�M%
�~=A�E2M����Dh�f��%X�W�>�tm��D�O�U���C\Kѐ��Bsto(Z>p��-�ҳM�gg�9'CO�=���v)}��I�������G�%��	��[T�v���f����ep���=eH��PG9�o�5�i�8�&\��#z�
^���=g&���P;���s2:?<Í�B�C=0)�>,Oe�8M��|zG"���kV�2H�A�X���J�c�7�ݴ�6��!S%`kB��'T"�f��	�/)�f �i�C��-�+ʀ�C/��ٛ�-��H^>��|�����e�k���4��x�zA�˺�V��(�
���d.�0~�E��+�K��VD7"��:��:�Qg��i4��8�[��˱�:n�d����뼀�_�止�S�b5Tȵ��)��C8�,�31�s��/�ލ���[O��6�*w&��O�@�,���¥��P"��!��?��,s/L6���Юiay*��$uu�q����D�����}������AvO�q\�3�:>(���2ْTԅ�SM�+�8Β���%)'�'5��X��8>��}^�SA��������yQ7Y���NHʩ�@s�I����Z\�ɸ#@�������ri�:?���I؝&��S�r׉Ó'SgJ9͈����p��IGx�ED7&�����廤:�n�[���e= #�w���y����E�hR��H�)�˥�{�����/���OLڞ��m_X�:D��_������褜`|�����f^�ܘLC?�"�3�N�ptF�/#�Y*�פ�����Ȏf��2R���5|3�½B^t���J�s{��8OaJ̈Z�򤤜��N�d��B��|~�K���Rsv	Re�sI9���p��'OJ����=R"���J��Q9��f8�f3��sR�7�ҁ�!~�2�՟RT�C�3��6��L,j~nݬ����Ƞ��z�9,��ڲ��"��Y��|_Z��r|��KF�e����rt��Km�zi���B,�������t[����Pߜn�)rO�Uq�gZ؜#t{RN�#,O��ϒ
��ߗT�&�W�
��FR�5��:!��MI��s�5��)�
3��|ί"����.M}7�vo��_�ݧ�V�p^8
�>)Wc5'�c\$弗Q[�)��MR���݂��GmX���s�K\�����V)�����<��]��-�a�\����Pn/�^��+�Wԧq��/07��������u���+�L���,uR�� l����X!���/g��+��^*�P�ϠX�A1MPp+�'y?�S�d ��9j�����Y#0s9�ČV�ٚ�R��|��4���n�}*����,p���������>�(|]x!��2̙���������X�̀����Ì�d��kQ��*�r�[�9�|��rr΀���X���G�����:���Au�Ɋi�#8�ӼPo
�H��S���tЁ��*��u|��_��Qx���5�]-Jxd�w�;+-�G#ܧ(��*�us4E��D�[��S�Mȭ�,v�Q>��=�-��a���vf}�D9�71Y��E�	�w	���?��Z��R^�I>]^<'���W��a��&�I�mZ1a��s�yV����]/�a�~8��!%���Qs��$�ɢQ�Ƨ�4DC7=8��/&۷��/4};�Ӓ0ң�m���`Pw�6W�e(Z#֎���x&�j�<l@��6̗V�OZ-AI�j�a��:�9��=�G�I�Z���M@�M �1�7�0��I	y4���ҝ�j+X:��$5ԯ�BΆB��$8����M)�&��;�	%�&8ps�	)L�L毥v��`{P��<�	��6`���8��)���^&lUj�s�
��l@�"MF�yh�:����Ԋf��~��s3������R7�>iz��/ôN(b;�$ݘ���)Z�KBt�L؜�s7 n�'��¥�얢^��u��cr�4�2m[��r����T�Jx���m��jt�F���'q��S�B�m��g/o���F��k�/�!3�:����msK돰��J9���ηML>;�t�����-�$�5,���1��jε4�,Z
���>]5��$��t�x�b�s��k�f��s��*�?���(�/�(��V��D�	�nҳ�-��ڳa��:�&c������1�܉:K?�3B+4}?C2��>`��9������hp���!�QgCE{�%H�O.�L2g�L�]!74O��e0j:�ur��qoR*v#:΃�K�[y3�l�e׼0�\�X�����DWw!Ί�1=��b��i���/	E�v@�E�3X�B�D�贏��ѝXWn���T�_G᝝(3�Q��#�;�6��g�F[�<�����9�GV7��X)A.կ��M2�Y>嗆�cj'�xy5/OO^:n��@ 7I��c}{�O�=/ۆ�n�S�n$�B��qU����G���_�&�l%#���J��f�A���M^t�����ߞQM��8���T,�T��5�DѨ��cd�r��l�F5ӽ/Uև�����ӕB�8`����]���/��yh�Nh�ş�y��O�#SC����\}����<�l뙖yIm�%%�f�����U�Vl[��֊M�B?�O��u�~��=��$Q�"�K��k���n�p�j� ��Kż�uջа�M���"��.A5��&��jS��r
m��B��j�r��D;�M �?9y;���߾�����Z���V��*F;�z5{aQPV�_r/���M"�=�UY(X�`4�u�x���O�x�)�G� �H��%�R��,��o��O�K���Z����'�m}̑���s�7% ����β��i+b��Pe��c-�R�1T�&Ə�LLY��
$�Öu�R?Y��.vp���:l֤)�C��4b�I���*�A�+�Pg����x������ٙL�y����u�=��s�����{���$�? �g xa2�� ��\"��w���v�z�� �a�L�!�Hg���aOs����,�fDpȭ��F���� �Hf!=���jh�0ߋ��{l{(�!r��I,g�-���$ڹx=�d��|W^C��[3=�b�[�H[cZS*R�ƫ0&U�n�ӄd�ЗkϾ�Rj��6�.w򻈀�8�H-�_�/��%�->�p��\jc:Y���D�T[R��ήR��d���6ܴ�.u(�aZ�.r���Z�F=L��/N�7�#�/�}!�<��v3�2a���lE�6�d`g�G���s�/Ê�M�ަD���p���Lr;��:<<��v��9 ��f�c+���f�>��/��8�a�����E./Cb��(U4wh� _nk����M��"A�ׯV�w�M:I��	�t7'�����������2/Հ9�?�4ɐ�EgzVQ�&.)�nB�c��U�;�%N�:��93u���uT@���+�t$��/�1sN�{���3�qdc�8�ؖ��b@�Mb��I��S��P�h`$;��&W1��&6��(ӐlQ�J�(�r��	7u��N��	ef����.���Oۍ���UO%ցf-V�k2;�h��Ɗ�b�rz��d�#��Kݖ_�Ђ�k�*&�7^�bJ����(q1���=�k)a���v�av� ������2ȑG
a�Zo���s+��4�+E~+���}iSϊ���}�\+��J �0�m���l�Y (����p�SC���s��:u��}��\5�U=i�q�؉��I��;���o�TH��"���f�X(픀Im0w�H>Xx����3~~�e(_J/�;�31��MA[D��W���}�R���[�P&M?;:+��N	�|L�>�@A�3}��%m�?��85�`��E�Rc�$�>���
����H=�LɈ�'�}g�\�#��<v�z�*�Kx�.WF�B˒��B�O�.��.`�DM�s�P~+����bil��V������-s���G.Iͩ˜���Lh뱓=%g�4��:{/� ��*��r7W�$���
����X�j"��T�a;��K�nsl�������"L~DN/���cS2a������4C��5&@����xw+�'��;�E;�k���.\W\�j�Orv����Au_r�i�[�m�
a���%ͮ�psXW�U�R���To'ڧ�Av)iv.j���W%\j%kl�;�O�	Nr�#DnOp������WҠS�\��gr5�ؓ���~FY����/�_�dp�����2˖���<e�$/��ȡ5D�R]��mT�]���μ��5=Dof�/��X��S��.���6ZO�f4���,C��v���h��Cb���É�S����}��lڊ� c꼐:lƊ՟�y�GM��)�D�"ɼ��1Iu��ޖXy�}���F��r!�������w,�l�O�V�[�]Jޯ'z۠�St%�	�?�^�cB���Nc�&��l�&%�����΢��t ����[���{��/��'FD+�EkC?|T�ih�A�F�(s�D��]	�� ����'m����2���{���^��Jp; x��n}蠅Fc �[�ةI���$�YEI��� ��@9-8p�z0
��{q�/Fϲ�I0e�d4�(	���8�:;]�FP�WW%f�껩���6�1��L��D�Abt<�x%��X�O[�V��k&��.�JH�_����_ӲC�\�˒���[){�Fgv�0;3`�={�z[�}J��Ε�{���=�f�ô���fIA �>o�~���F,����yW�w�)���]}!�'ݖ7M_����ױ�B�E�.
��M���F���C�ű��Hs_���˱��T\�P]��������Q-�}$�I��ț���7juiw#>��c��ٱ���w�f��.�k��/8`�O��N�/ĕR|f�p���ğ���i��>�~z�3��U���F�s��eV���9E���n"���ǉ�Eg�ˑJu�q�K���y�?�b;iT���uC�8��Iu���>�7�±4�	������a�R*VyhK'բ
᠖RqZ�qt�(z�X8���.d}�k�X_t�-{���4�A���fR�f�qf�Kݕ~��t�V|��Y�sq���L4��F�R�T�U�F�(y�r9��<4�lU��8MiP/}�ٜ�A3�<�X���R*F���v�1�_��Rɯ�:$��hМ�&5hNN�zhN6�4#�s��M�<�lS쐙�X1�_�Bc�{V$�Ѡ����Ӥ��fR�f�qm;�"�2�b���܈)|~u{0��Ww��Ѡ����Ӥ��fR���#�bC�8��R����C��eEh���]t�[��[�-`�fJ<��P7eC��>+uK��sM����������s����t�=���\�"��\{>gN�ek���p���DR��l\{�y���-3מ�����|�����s=&3מ;�����Y����s}*uȵ�����2s��������\{�j��^��k���?�_�̵�-���ݙ������P�\{Nl��^��k��?��g��s������\{�i~\�
@4�SԲ�u����@�\M����C󜃈kb�<	��m-D��x]BYEF�+@�CQbC]�j���n�]���C�z��OD��QK�S��8���1�נ�E�w�ė���4��_��U�dr,y$�{U�ּ�|-����A�F��M�bm,�-��k	�Y��fa1�I�T6�]�[Q���+ɗE2 ���wD݉2�Q�	v>�����c[�烙U���a���?3f[���A�zU�����Fj8���<�Q]Râ�Y�\^uvb��Ύh�̣ٙ:;�yTg�.����Q��+�z����h�0Ai��0�kY��55\��Kcj���=�ἓ�7���sV^���v��N�>�n��gY�!K�:1�m�B�ر���5�s��N}�&02������3��H��|)90���R���T����Y�a��2�](���xt~rc�w|��u�%�kZܒ}��!$�8�����3�o�&d�hx��"Fs�֍`�!���Ӊ�����}.�5/t?�qt(�I'�I$5k�r���ȬWs�A�ч5��N���J}X����B����\(s.��euW�y[�O��=|j�Du��l�Y�O��I-�%�G������pH��}ا�x��{��*�7�b�7`e��6L��s�MZ�a�>�"���ݽz��<�*����?j�mj�W�ϱZ`��)tQ���]��ݡ�E=IQOJe��i����PW�C�+�^�O\�	�`B--ޮ�`��L�<'C�&���qn���B�:f����x3֫o@�[����AJ�H7٦�k�2�4�Am$P��o���������(�m6��S�|:#U�R�	�����(X�����\K]\[]2�1�|Y�����cMЁ�CL,\�,jT�j-0�^v��?���)�֏�8S� F.`+�+�,�U����Z��3�jU,�n����d��2��p��t�x����E�Y�=�E�T�¸�jl*U[��d�%���*F5�!�!���O��ꈣ2Rׯ)#rL�Zk��S���|��%Ɵ"2~LdD�������u�K�\�R����K�(�$7J�!�2�&�Xj{ҭRH��=F�UYЦ��R��(6#�L�L�����|�s����w'0��@�rB��ж�[1>3_���^�V*v��fע�Lz'`UD�S��(��2̃D>�TGЏ�m-����N����錧Ka�[C�=��.��j�ڟ�H���{J������2.kڬ(852@���x���;�4H�@�K]X��*�C 2�/IJ�����2��@�6��Nx/��"Jۻ.4��9:��"@kVh(�֍�3���Є�&�Lue��	��$sڠ��Sϕ�)w%�vԅm��� q)B+���ru�VS�~�����zT������XE9�V��pߋW|Ƶb4����/��>���'�7޼�_i��Җ�+B>B��gp'��B5���� '�aR��Qwd1#����]�Aw�'�t��8�^M,����A_|�.����V�K�&�zgi��*��=J���
P>�U��Vɨ��m������в�}-b�)���Z%^j�u(��G�^�z-޷Q�z��re�0�M	(
���o	E�N�6{�{���(<Fd�<ⶋ�^���eԬɛ#�pXŮ�O����%��!Y��t���@�L*����15v�j�u�>6v�I��R*7�����U�s�Z�W��u��~ꝎՈD�i�]P�J�(�l�f%l�k���a@�/��]dy�����!��� �=� �>%�b���^N�Ġ�@����w�먣�rx��1R{ୁ����L����N��=�*����uzM@�޾]�g��4<)yS��̂��տ��VN��M(�K�Q�~�֟F��=����kU\rA����9!c"���K�i_��4\�^k�
��Y1ʵ�����U��@�uu�
��~�.&.?,�|�(�]cu*���_�J�D�@�C�u���o�~��j�=�;Hï�x��F/g�����b!���K�+��ï�>��8TC�I-##���9-�u��Q�_D(��+ud��ۍ)p�{������0�v��������N���[h��2z/#l'�O�r�Z�b��K���oZ�5��}]�!�����W�Z�[�M�U�_U{���R�\ZRU	��K*����̃B��O%�i �l�D�ɟ`�����S��T�9JK4�����qjb���H���l��HR9�k�p�K^ĭ�G��{[�f���c��F�z��{ɧ�ԫ�Ƌ��@�{NWG��T��]� ���%�nm�����7�Рe�XIxRu�#V^
L�2��e�Bۓ��C%�@��Ђ���S0דՒJv�@Qx ��2���)��v����u�o������\�gI.ܧ�l�����'����s�ހ;o9���4��@�)'@�gB�"w�N�jB@U�ֵ����nP��4PF��&��ß�g�D�͈��,W�mP�}�%+�hɱA�Ԁ��J#�������/"+g������;i(��	XAQ�D
wR�o�t���X�|.��QG�zw���ݜj����F ���#��G�������^�`e�\悵��W�o9��/�z��ʥ�7�K|�ƫH�媁�\�u�ivi8�fЋ��)�!LgY�r��q�jw�b%���O-:C�W�u�q��P�0�������� �l�S$مV
�r��A��jE�#��,z '��jy��N��jA�P��=��L�%�>��*� �X�Q@$���)v��^�f���=Z~.�����z��*�R�S�u'E I�Y�HT�Ӱ��]�!���t�Y�i�aIW�Cdl��9�p<R��9σ]?G�I�vwF�J�,�R���z���W` ��7�C�����nI[����ѿ������{����b-|����2x��~"�7s�$Rѐ,b��wI0\����*��M�C'OV��D���v7���J���v��T�I%�,R�S<�}�D�|�F�R�M��_@�JC۱�R$�ydv�m����~��?6P��><����.��c��ޠ��?��T"��Px��b�������"l���Y��4��$��Pt^�@t�������Dj�ئ콊�8�T��zA��n��O�
�"=���`���q�ysV�5x����$��[�X�O�r*�"�؋.�<Za&�}m�-V�MOn+]�&%ptM����d��1�;����H��B��1˷'�I�W '����n�
�t l%F�>�X6��	�����O���d3:,������0V���z����X��e砶Z�;�Y.�.f��C��O��/pT�_E��,c
IL��v�
���?�� � ~�-���
p�+=�p�fJ��PQ��s����>3����"	�h2�#c �u� 4bW��	�gZK_� z�dBg�K�K`gF������	��&z�2x3�x6�;OJ��nD�� x�@�}	u�C1����H�}�юµi�e���*)���f���A�x���)Fn�cL�Y�$�w�G	:�|�|����<�:Q��|T�:�����$��g"�q��>229�ь�4lX��������Oވ�x?Co-�v�ǛQhV!�o��Cf�DW�芀ԂW<O)�f�������u���)(�C�ٌ^�j� �i$ݞ+afs"(iQ#�e۪�y<�si�]P�-��q��?G1��o�=�&�a�����rP|�O CAQ�2gb��q�&[$Z}(p��_�c,
_������DZ\�+�ΤV�qsfl�l�	��21Ny��� �j�Zr���G�Q��V��`�*��`�FzeN'�L�6�Պ*ʉ<Lc���{��9�>�G��_�׳*{�~��")QC�Q��M��ֻޫQ?��E�����ӽ���0;<���Ձ���X�WA�����S�Zi9��K֝n]Y�`��A���A8�a�u#Q"D�*I-���_��RU`�_�0H������@�	,0���!�� �*�e���]����*��SJ�hWD��u=AkNs�҂h��jǟ�ga�>Շ#���J|7��u��@9��O��pT�Wf����Xkt6����o��`i>[=kƪ�:�Q�}:K�x7Y�v%���9s��J�$è��F2�ַb��E�V�����#t�4�)�&��-H������������ �Wc�@Ӈ�h��Y�T�ڭ�u�V��(��gZ8�Rz��B܅�IP�$(�Ot�`���N���FJj��U�7At^jI�|
�N�����э��w&Ҋ��M�kIڞ2�|jK��t�ۓ��r�I�Hi�+<��5T2o[��]҈ձ+rd��
�X
�-S��?�C3;+ �/���jD'�����u�_ě�9JYb�9%�%��jG�S�&r�~%=W��mđ0[�ء�&js�d��'��:��j�Ō�C]��m����llM��W�Q�A������bh6/�<�#���|���Aj�q�CѢ�s0A��->���i�Ѧ�U��X�\�c[-d�[
�2���D�2�1�2����^�_��,��T2$���X�Y
Ϲ�v��Wi��	� ��$p�<NP͑�+A�ݪ���MB�=������G�c^����;�ؼ���ɜ؉�!$0��U�AAU�P!'���vb;�?b��׎�~���o:�ҵ[���P[+�U�uHsl-e����h�n�b]ʘ���R�i �>_=W�����7�t��ի��s��y��<�y�sι�6���r�4�������:`��&΀��߯#���H�>n+�{p�s�esy�m{�-

�S1���m��L����i3���Z���Y�~�v��U5���T�~hʯ��U�X8�S��b���Pq;!���L���)7��G��|�Hf2�6�7���,rs'�L2B
�#��9�K~*[�j�UO`nӾ7~�J����!����F-hn�q�]��A���T�<��SQ2�l�?�;�� ����5ȒO��T��S��
d�r,;��ŦD>)@J|�ܐ���}�M�4c rE*��`_J�;��?�
��;o��{G�.���\*�'|�R���W��+�G-��������Ŀ�H5�ʽ~����UJ}����Y���7��"���E��?uD�2���ϹF��a��4 �j���T�ŎP���DR��O�+�0�/����t'}���ÀO9�x�x�(�	:�1P1բo�7U��$���ێ!�~�ܛ���[�ki�/���T ;�=�_*�)y0�+�-�slsE�+��i�c��}�@�}�H�;}�<�
d�?>����}J^Kr�y>U7�{>���J%�+�e2H��N&-%.Ⱦ��<�ڻ29����C�}
�G}JN���o��Ril�ggG*J���\�
�M_�nN���+x)���)�>%7���"�L��A�H����T _9�2y�)MEɭ��ͦi�e�B*=y�g�<�LN�]�|*v^�]��iA\vIZ���L�	il$H�^��:Nۓ��ԡ*�*�N��X�
��
�s�"/����Rɓ2tx�:�f�i�3܊���P���<U�ݩ��'l�'�ƨV:���,��1�KP��I�.��r�s�͠�	��?�:��C&�������h�9�H��Y�I$ȏL�ɢ �Ā\�k���F�)����ǣ�+�纋��X�t�t�+<q�{���î�:���$`s��:M�������<ḎE�Ʋ�H��e�Q�����שR\	����T �}J��
|��9,��a�Q��i���s�T����"�J�5���āl���b�@�����a� �2������T�Sr���	B ��px�I��u����t��]�}�7�������(�8䃼�H�i��,}�)GI�*�3?��Y	%n�	���7���]k�r)�8��XQ��b�g����y����
~�Q�8J��梿IL~���+���0 Z����%˸K<y ��ؓmLp�p
h5�WΓ0���țN���y��r?Uڝ��~�$П s+j���}��B��a<k�a�Α���*�Rb���Sk�r�/���@����*��Ǐv"�� Z�Y6-�>��\Z>��ub/�B;��H��]���a���H�UO�TM�d�vQ#=��p��N�X��d��U��P�|��tH�fV��;�SQr��?ȗ}��T�Or>4ܬ����]�~=�ւ��7$ә�>UO�X{=k��:�3T 	�I?��r���`�ϕ�CEW�I����C��--8��{�՟��cʀi��^��a>C4ss�㮨�/�.����V��צS�f��b��o%�ꮵ�L���"�sdR��}1���Jz���]�թ���/�#)�)��#M�	��^�]�����q��N��vfvz5�����`�:s��N�x�h~�Z������e:�3x=��ڻ��u;�V�q�3��|���zM��A�^�g8C��O�|��b�[t�v��E�ba��m���z:�w�-�B�Ù��]�?n/�2f�?��1�'�����4�j����o��\)�7�.���|�������[Aum�=oq㧝�����w�Zk��O��"�k�KD�K��*�.���~�뷈.�ݽgn������'�30]�>ڪ%D����c_�a,��=�	-!���3�vb���;y2�� '��Q{I�^��ÿNAj��(�5�ғܿb����+�<	��V�I�N0?�`u�8��k��:�[��q��/����M�x;�����HFۧ���ݐ_1�@2�Pf}�j��~��=������㾙���d�A;���E��-��⳼�+5�*`S�u����Wi�<T���˺�|�)���;G�?Ǔ���`����y���r���e�i}��0��p*W��k��-��&笝�;��R�޽��t����s��s�_��n�Y���ν{�h�S(x�v�� ���g�-R~�r_��ܯ�_6p𰌌�:VC~��kb*ay/��nN���Q�[9��|� ��!7w}�#H7��?Ip���4��	"�Dt'����>��W|���Z<��l[�̷1Ӽ���-��7�'�Nn��%�������B�1��	��!�G�4=����s����`��ة�SK��j��fG9Y���4�ƃ����;�65Ĩ����|�	��6T�2暽�ת]�^���]��ʗ����]��ɮ_Hf�?Hl��.6�EȮ��\�+�>$v=o���y`�î?jv}������Z��5��m��(���Į�_��:��L�g/�����<q�'�����z�c�~3t�:�o��\�Q�g�Oq�&h�b���g����A����$�E2�V��e1����/��_���n���M?k�]���m�Q������|0�g������:v�C6e=m�z���Ȯ?ϫA��>�X(cw�_�t��k
��;���0��K$ۋ)����������K�Y��#��XyY��W��j>�}�V�ݿ���E��l��u�'��U���ת]�^���u�>�uˢeݲ�X�,Z�-��uˢe�U�{�)�f���(ȧ��`��L��̛[[6��~$�V�z�����R~��w�_�#�}��:�Z紵�V�6��&���D�>~�^����I*�	=?�$�|��*?�@���w��(�.�Љ�H� g�����	��b�ZU����*�n���馣��nF��ڪ@O�(�I��B�,��� ��P����h�v O�b+�Cg_��du5�F��`y��1y�^��tV��e���u}�]��һ�kP�q� %�\�����q;P<�h��j��_��3�)_}���sa��_�_3p��C���嫗'wA^� u�y�ʟ2t���eǸC=�W��]�Cp���8u�����h��}�����-����[�쥏b��<�=螶1�6̿�FR[�N��s��ZS\�m��ix3���È��(N\�!�qf��	��t��[E��YͲ���}��K>��O�n��x�c��?�i�f��� ��S��@m;��a�����Rꄪ	���rr�2�d��{oBÇ�RA�.�`"��m&�9p������7ȝ�Etb�=����� y��Ӷ�o7�;b�Mf�i�����KQ���
$�o��v�����W7���(=�0��I�-0%=�̟mf��Qz�#�� l��"t�}7�L���q,T�ю�r�+�1`�����.���m�F�1~ �2/@d'�)���*C�H:yj��_YF�v~�AրU�$�̣n��2X@O+��{3�Hn�~�#��k�2
���������z�� ����t��rP�AV��p���P_Lٗ�r�����$��,l6�3��&���Yz;d�[������2�7:��ufV%�Pv�/'�+C�-ܻ�c6i>y��@Fikrӧϧm�R19�쌂<�����b�F����@�ct�,zv�_j�Z?��ݩ��-��I�>��c{�mG:&ۙ�!I:�bF ���G�sԚ�7F��PX|��ED�F�h��R���o��e����.�y�cP?tX��f�أ))�X	��fA�����9o��m�tE1��Xgjy��H��:�����G�tV=�����Ɨ�<��.�5
� ��K�|���5Ui1~��r<lࡾ��N��'�~���WP��&��uLn�p7'j+�� �vPE}]��EκRo�i2�.��g��"5�"���Y���������J��b����Y��\�}Z�Z�ƃ���Z�⏘�2���xX�mFꐞ�//:J͊�� hM�9r��u),���x�xl��z�-��؂�kS�Ɯ}lK�6(�+J�<�8��-�<o{�lF���{��׍�����j�ZP�0��g��#:��Q���^�+��|E�d�d��O�r�V�<��x:�k���9lmuǌA�ǔPy�+���
�����E������9�yA��MC���$�g��>���qz'��ö�_��6wT�˪'4��v����7�1�@�����i�U��D����fn�fl��X�� ��Q@��&�c	��|'��l���1���9��
d8`�a�����J�����1tjL�30~x�14_M�X/�i;���G�'T�3l�B_Uނ�]�`ī����i��F��Ɩ˵6'��D���y���	���m�J���p;���O��h1��1�6�h�\��V�n6�A���>MXW��F����V��)�m{Q�~o��{��c��L[z����rP�،^�d;-�AaxN��Q�cTY���ʑ6�����F�B9�6�f��v�e��?PS���a֦��T	�p��簁��0���S~��n�3�(�M�X��r)O.��.m[���UΜt������c�#�,�:`ߚ�6{�Z6�����H���h��5�#)�,��.�SH�-5j�qQ�Y�I)>���<PC�G��{t!����U\�5K�C�,�	�w㦟���L�OȘ.��o�Z<��� ��$���G,F�-��Z�4$/�e2l5ߢ�-�t��-������.Y��t��b�!��3���\��7 ��;8zc�t��rw��F����!u�'���ԛ/v��ݘ~��ϸc�7x�Д��(�/[�1�3��S��n�/����m���JЮ�P��
_'5�Ѣd�sP2ocD���4��o7"��U�u�x�L��3�W�a���ļ̛k�l���?n2,1��!��� �'`���M+JCf#y����J�J�1?�dsd-|Y&�����FD]M--d����i�9�>��1���GͿ�D��י��j��T�#	�Q�pZ*���l6��J��R��k��͊w�lk���RJ^Շ|u��MM���5�����6��7c�(����P�������d����7KQ�(Ym�XQ�X��g���^�iB�\S�:>vԔ����ֻ]� 7�1}����V��j6ZG�z�͏j��hM?k�Z�ɚ�m[	/�4�Y�������賻Fky7:�� �;Bc�^��0�ȰG��.�M&�4�J���Q��㡽�����48V[�z����i1o��	�4"�Ƚ�'S#ml�ˡ��X_��\J�M٬6��dM���g�d��Vʆ靼��MP.ڂ��`92k]�3~]Le�;�]��)�����w��Й��s�XƔd���v�E��ů1�;4k}V~^1R����Ϝf9'��i~�o62o~`��3�`j�t���-i1����Ĝ�7`2G�g:�Q���3k�)����'d���<�O��SE˫�,"����7E����� �P�w�X͛�x.U.�61wq��Rg~lohO� v�J-<� �9a�:��h��n��c4�*��q�\�b�a�tOj7/WW�N�Hek�F�֭:1���]��#h~+M�8AZy�-�&�Yy�y�w�"p�!���~�3r��"��m�9C�����ή	��(��6x���T�-E��8݆H��~C`�<]K��|���Q��4CU����
M��C���w��Z��z�|c�w��Q��;��M���`�u���B��|�Fn4$���X��`���������k_�rO[G�u��ǻ�VʣVAs`���V�'�G+�М ��ec��FCP,�G���}w�m�;�Q�K�c4D:`N)|�%��Dss�OP��]���:�0�I��^�Y��Q)�&���G�i�}�	A[(|�P�	�R�nQV�)I)�7�)�R��b�T�������M�F�����S�S��E��ЪV֔m�Z*��k�_m�T;7����ʻ}��m�7X^\��E�e��-�V˟�\=��ҕF��kaC���w�p+�sN݀�A���e��p�-(�>=��7�aJ��-�U�98F��#�f�w̼�K4k��9���_(>	�y�h��!K�mE74d���q�6f{i:-�=��4����`s��
*�T���E�����G���W����a�"X#�U�0d1��yXh �ζΎ �	��p�F�Ö������̿�4��c8=i��>ӄ� O����y3�@�� Ϛ�L�)W��1�+Ш�M���y^�V���>�ϓ���AІ�Ƌ�]0����ˣ|x���^N�~=��7V�ٶ4k,S��l��'Ö>�=W=� �ߍH�mY3�w#gwϹ���C��׹�1�3ˑ���*�����-�_B���W�4�� 5�o7Cyj9�l�A'����e��E[��H!�=������FT���Y@��lC��I��Z�si�G+A�pm�ڏ'l�p#Z:c�KcD'�= �C6V�t�Y"�
�&nM�fl�*��&��������v�c´��K3;�$��t�@�H@A�a�COA�ټ�a�3���l SQ�ϰn��+�*��L���o+o��=T�?`� �u���7�ޭS?5��9��(�B��
�6j~i��#4�	�������[*�֡�jd����H�}蔙� �M��N���$�7�B�xT̯�@
L�_ՙ�q��]��¬�)Y_�,�_j��D��vk6�֩�
h��xc���;����k��rsOn1jD#u�3B�b�WB!@H �����a�@���ĉjiA�糈�����=��"�OD�(2
8 u@^���u>;w"������|?��s��g���Z{�����+�
J{�#�4���vT��N	6sc��m�fNcx�ɭFy&q�G�x�L�����q��L���1�Й�W�E���Q`���%px,y�e�)
Q�#�j,��S6 ���8���V�N�/ +���B9�R -\���b����qI�e^�m�P�A�h2���d����g}I��ʀ�Ii�"�G�S���k��֘����C����!��-2��q1�O�����w��e���Oa �^7�Z~udI^�-'�/)�Z����W��1��M���1Kj����=�\it^��9���JE�U�Y�|�:k&�f^jPß�\oJ_{y�3�_aM{��9,�]�a[X�eSL>��/�Or>�ڵ�i�5N1�c�6Y��R�!�O%'�b��tƘ��e^\M�oIX�3��׭N�tSg��z8��O����r�6E�����>���4�Lz�]&Sf+��;X��rV�kc�m>B��_O��5��;=�ce�^S�Cqھ�~�A�����l6���1s1^{l�����39զxN�S�kR���SƯ�=����E���M&+V�P�V��o�jzr��2Y1=��D�}v�y&üB)�P�F�c�E����٦��ѯ����YF�:��yD���޷�iDF3=助6�_K�[}����9�Y���k-3%��@.�}k��U�C���ì�PO�rl�Z����h<ӳ��ޓ�#��x�Y�i�����5��R�?�LC��	�9F������b26��Ϸ. �)�TpN�dYÔ��yI�q��lW�y�i%��|;�Ɖ�l�ʟ�>'������(�s��l����h�P�w�kVP����d�̆D�Z%T���h���:��ޑ�[��L�V)��"~���΀:eu�	*��|�z�ݥ'|��fM��r ������~�]X�T:�X_?�P=�i&��_kB��yK���D��MC}	���ӌ���Q��u$�$K�����%�ӛ��?�F���.ZY"囔�~��䧊鋈���.!<.N�u�o"K�2��RL�&����}-�#uF��}:R���;�}l�����	����ywH-���i�w�˫�F��_���Y��i:B���즑g?����E����|�d(a�T�/Ør���#� ��':������K�}_��k���SO�:���%�ƐB1L��J�O�Ʈ�x���6۸�r+�i�ޚ����A2x*L�KgX��鷋�|�
�����0�q���Y䪪cs�������'5��h�l�0��7'\�F(��ɣ�>��C��V�ʾߵ��e�$x���<Yi��j+j��I�I����ڷ�k�J�a�\�M��k��ԀoE���7"B�=.^��<���z #�U����H�"���b�$��$����9S�z��7?yY���\L��ט�4�ʿ��{1�'��S5p�Tm5mAMF�tؼ��XV|��߁�/
y�&�]��q35�������7"�(�w���
�e�/� ��w_���bZ�"���+8�Ŏ�/���&�WD\�����`9��k�1q1��剋lC7�j6e��'ng#�e��Pύ�ن���`Kc�&ïq�j�k��%�x���ZO���F[��IN^�4�&�3Hp7�\MYm�վ�S�~���y��ݖ�$�<d����b�6ؾ�s�<ҙFn�2+j�黍�U���]϶{l������N9�$[��"���?�θe>��Y��]|֍H�m�������w��kfr�N*U�{UR���λ4����5��}��Ք�j
�#r��z���O�A�yәV����ei.���9��?⫭�lw��*������_'�+b�A�@�VXXl}%91dhG:=���ۣc5��]l-���B�8�$�y�%���t��,�k���g�m1�߭�=����I��pu���F�7����]�w�57�֜�U�R�鏫�#���ˊ,��
�S���\g��([�i|YW�Qln����9�r��)U$�5�u�L�8��p�)��'k������!fD���X�_j��5U��'*�T!Cr&{������W�)�g���X�x�H�O���x))k��&J����RѩO4�߿��cEh�a-���(JP���PhZ�J+N���VZGCS��Uj���k�Y �Zp�r�	e�ɧ&�)H4�`з�����{�����|������9P���oQX��.��]
w��ޏi�:�G+.��|�U��z�������:n��j0��<�[g����Yd)�:�u��d��(jW��qyU�c�(7����DY)�@�t+�&ZbM�ӡ@�t���2st�@�~*M���{0�l�nјi�7�~b��'9%���o�~�ݨ���"����j=�BNVY�ou����:�"%�fia,;V7&$"
���461��1V��~��D�A4.&�����XJ�(���̪��6!��d����v�f�+XT�o	�\:"�m�R�鞉>=�k}���R�����y1��L	4X�C0����Aj�TǏk�s�"އ��A��p�	mm4] ߏZB�(���0��o#M�[�
J؆̯��'�O^}���s*�Y��(7y�N��K���R�,O��W���q�-N�^�m��=-;si�v=������	J��y��ܯ/:�<�c�Q��ԙx�U��Sv�k�h��#k���x\�P�)�|�j�#~�y�|���׃����m���p��H�H��))��i�4�K�t������G���F^Dq���X�o�X*�Lng��*�B�l��Q|��C��X-�1�.V��\���M�'�/�`=X���U.�y���N7��X�)���+ٞ���U��g��Ռqd���;~���4���V��J\O�9t
�����Mk��T��9Z���'*>v4�pv��E2h��k�I�j΋ƹ"�m�Z���[@c�9V@�̢&|��i1�XOR�ݨ�2��Z�i�#;j��{�����r�l�!&c5�F��բ�uC�����&���=�?�N�@�9����÷Np}�=G4i���&gŋ���Lj��Ph��&�l�����X���4�MF�x�|wZZ$Ţq���b�ufj�Ѧ�[c�g�ͩM���>U����ZO�~W�7��M��.���Z$��j�=BJ|�]�+�[F@Ei��R�!�B.ObI����r93��SDr)�!�B�%=b(��/U.��o��i�t?{S=t0�Ƞ?Ǌ=.5�:���Wg�+���D���:�f����K�M'��^T�^�F};�������
8u� ���r��hovR�����k+�K�8�9��α���9�u���T���+���/wv7�ܶ3���5��,"͊�C�=��v�k��5]y���#�w� ���z�E`��::E�թ���GOr�S�s>�n9�����)�\N���n��_+��:3ܩ	�U���X��G�M�j�N]mtZ�4�n+\!7���9�v���Z�@b�X�BMP���Uλ+@�"�Es޺�)7���[�S�����r�PɀQX]�{C-���iS��2�`j�>y�ag�s��誘9$x!��~����Ӂ{�{{9��#�C�4���1��G=KC��:�|�9^�W9��9�,q��󾧰!i�)�
�����:���K'�u
dZ������S���-�S��;�*L��V^D1��T�R�����U\ǥ�p��ꉚ�k�9Y%W<��F���Jpr�5�1��=l���?���R�k�,��I�&Z�$�h���|�w�w�w��O�;��?��{�v�>IG������s8~
��nP�ݮ�y���P:�P�M�;�sa*f�l���f�~�ȹ���Mp:|�O�(�V�Z���.�'s��6��ͥ�~;��i�3�	��	����zx�?��5�m�.�y�j=���Dx8�1�d
_'�<��Vu���!0>���������[���K�)|n�o�W�+�B:2��3�	�hx���A�r�:�o�(8���	b���G�1�\ ���t���7��p|��Cx:<v���,�p*yNźH�jJ���J_ )������G�����g�:�~�7�?���K�9x��4�}x<f�U� �S �;@�'��?���
`���m����{��p.�g�=p'���up9|.�����O���H�5+�j4d��C�Fp�����?��]p�%�����p-|�|�G�?�����pl�S`��y#}ɶ�U���?��	�·��_�u��n�[�;N�����ED�O����0j����f�%�FÑ�8��O�'��Nx0�o����3���+)ۥ?]��^A�y�Y�L�2�H�t��nA��,�R���-�A�5h[5�����~x����n�W��u4ݻp|�
����?�g�c�Ѱ�Lɶ2�U�@f��2��Z�)I��?������+x�N���'�C��W��7BOx:<	v�A���`#���P���?|>
�{�<x+�^w���p|���`2v<s,�Y_˞}����T�͓�j�E[:*��i��-��ƱRn�3�p'|��o�����K�O���0�!��4��m�&�QP���([-B�В!$a-�M�В!$a-"$>��!	Ch��0��!	ChII�%=$���TԞ��
�CKj�M-�H!��!	=���$�В��CKzHB-�!	=���$�В��CK�q|	�	^��;~�Z�4j��z'��'p$,���%�I�0|��?��r��=p�7�up%|� ���<�
��G۵�j�
�5;�B��t-F�ђa$^-F�ђa$^-F�ђa$^-F�ђ��|Y�<��],þ=* �^ˠ�1�#�=��o�3�n�~߁o�e�yx��'<���b� ��Q
Ϗr����|>�;�<8^����g������0�&��	O���k�A$^mD�i�� /�6"�h� /�6"�h� /�6"�h� /�6"�h� /�6"�h�T$^*�0���6LE�IХ�O6vG��p0����x�N�_�O�{p#\W��a/
���tx<��gYeNF&��)�d�9)�L9'#��i��h�dZb2�0�rNFJ�x�a �@�x�a �@�x�a ���6LB�%���xRܪ�Ih�$$^�0	��d�=E� ^���{��p.�g�=p'���up9|.������0i�_έN9O�}��PX
������ ��k�+��Q�~7�5N9/�*�§p|,<f9��Q�:���L[��g� ���ͭ����#p%�����(��p�·����d��X��J�|�h�i��0_�Ci��,��k鈋H�(X�vl�=0�{� ����Y�+��������R��h�T�I*Z�o�n��*�M\����< ���(��8>��Y}2uo|΂�P�����(&-^�!��gހ/s~1��t�����`t�ڟ�a��95m#|�?=�Iե�v&��z��nͤ<3)�,$[�2��i�}�r�Y���Է{ɞ|��z:
]K���N��y�<ْA}���ˠ���vh��Yr{:�FҐ�!�;��[��#ߠG{�����e�S�y)�-A,� K*�[�'����78����=GV�W���Y���{��LE�n�C�0N���R���p��$�H�dj��[x.t�
g8}��/���9N�]�u�'<�:;��]x�4�}��������]��!��U�|>�wdׯ�,�o�W�n���5��Y�/A��s�Ư���P#��P�}� ����M�^@�<��4��ǯ����&xu5ّ���^�G�<��톛�:�_��Wg���,���x2v�3��A�ݱ��|���]K�jbH*���﷬�{'�\W�W�	���a6ԯ	N����t�z)HT�_-O�/��p3\Orڲl���p!�.w<�=`wǣ;±9���a��5�Y ��]!�a+|�k���5Τt_?�������w��u��k�6m'��Diw������`�s�;�g�V�?� ΃+��z��,�]b��Zpu|>5��5EӜ�C�[`٘?�oC�$�h��R�x���q<�֣�{h�4�g����1�]��<֬�0��0�ַaPKowFm��.f?���uP�?�c�L�(�=>� �I:Q�\|FmX�B@�+�	  GH��~P�N�d�$�pѸ��*�x�x�+j\QqA��z�x�O�c��E�f����?��dB�ɧꛞ�����]��w�Ϭ�H灕`)8| \���n �!0g�=���f~)�	p}�F�i�f�Rұ[�1�}�'�&p
�Bp"8
\n����L�|+�<~(��%�����DMJ�9|�ܪuI��.}ۢ,ǂc#��Y�A�P��y����$�����%�����Ƅ�vO�]���I�%����h� ���6���H����Az��t�^/y-x%�#�<�i�ާ��B���z�֛Az܅�s�r�u�jM<x���� _f�d��	N�%��"d+8u�,Ђ[@o쇐�Y�@�iC�^��o�o��Xk�xj�<pk�o_7��P��;��ԚZ�\>�� �R�Δ���'�����[�dEB����/�� �-�F���2��?؛��h>ؤ�7�U����4��Zk��Z2�T�h�q��ں9i�if��zқ� ��+� ��ޠ��5�'��� �U��GU= �.��	(�1A}"�Z/K�'���`�V�k�h���V:-g"t��h��������Z�K�Mj���B_�x��"�csv.a�o�Cج�^dA�ԭ��?w0m|��$�r���՟W�b3kIEa��Lև��F�	�&@Vu�y
Ǵ�'�y����x���pd�x� ��f�p9���߁�!f3��7Yk@���i=�nQ�R�}5X�Ɓ'��c#�ސ�߲u�	�#l�����1�w��0����O��;���)�b6>�$T�V�&�HM8�	��	Wjلy�	cJτң�s�VY���E�
|��������Ke�ŬG; ��$g�2X��G��
�p!�<�|6�z�٥l��&�C�=�L��l��lO`s�~(��ld�����gZ�F�'�S��j>Ӻ_�n�h�h�{`n�[�| ����)s>x9�Nm�L������{ �B��)����a�N��k����"���
��Ƅۑ�K�,]��O-k�G@~���hSo���c��lu�Ɓ���!�+�}p<$�Yp;���3�^�\6CQ���uw�W�����(�|��Qpx=[~��������'�+�?�������;��z�pӑ���f��/�M��J�.p9x5�x3d~)����� �..<��h�����l��l�?� ����4������諗o3{�� ��i*jٚ ��m�@z7N��'\�y�j�0	lfG|9����V(R������K�C�b�lu^���@�����7���H�{�V����*��iG7@ �?�
��Rak"�X�@c��٘V_u2���%}�HW��m�A�K�dqq��i���̲�l*�1�|�ØM���k��gl��8�j��oQ��i�Z���LOF�a6�
�$[��`�TXo/����}��¼n��������y��������dl�"�PoC��3	u<	�/	s�$��I�q�0�I��od��yZ�9�Y�/@,��^����oC�F�Hv��OA�ҧ�h~wH6[�T�B�Z�K���,L��a �׀}�����f'�C�g�*���L�x��j5��۟�궗���F��Z`�z���^o	�u��-Z]�^҈9�#����/�牲Y���l�������K� ��z%��=	�`�����,�v���(�d�S��2��x�7����Np8�.����c��?�^����L�f�&e�Լ���g���*� ��>^��tѤ78��H�l�2뎷��,� ��5L�@#���8��. �W�+��l̶���I�������"8�v&x����N��+p=������v�)_�lVG��z�Il=h8\�����6��Rt ��9lm��=W�9�u�np�閜�T���dq{�A`?�n��^Za��)`��b'B!��ӻ�p��5��q ���`6���e�6
H��� �lU��Y9�ׂ.���ɹ\��J��1m!�=��ʬ�aZ�����_�u(���a+So0��Z����,�/.���8�i�R؊-�eW�h��}�G+T���Bf�:���>6�e�{�����>HB��ʊ��@[�d��$�Qz/�-h�V(F��H�B��YL���b��@Z�H`��g�1k�Jp������<��� I�z/��%������5�AZ����ogO�X5�oX0�&�M��&�� �{�f��)�n�п�k��붅���e";�0,ǃ��;����S�~�=e�
��(�f��^�Z�St%[����Z�w��;�<�e���5Gisk�~��`O6v��l3�M ��?����Jo�����S��A��"%��׀� ��L�q��Z�t����o���^w��f��rx�֏��$g���i ����.УO��T�zQ}^�~Ƥ�^X��q/�K�opt��ULoCR�#F��m�6�Ϗ�&}�.���iv��HR�[w׬>����J�3�JZGN�Tɤ�̐�VO0���jZG3�HwHEw�ٱ\f��>�����a6�d�tӅ6�?���~p�1�!���na���0��	�Ŭa���ټ����f�^f���s��x0������c�b�!�6�T�2�KϦ���j{���lh�eڃ���j�A+{fm��%I �)��5��f]���=��m����Y�1I͞k{�Y���m�5�;�X�zf�K�뫘-�f�K�q���mL븙i���C@Z����9�TM��ƻ19�����j��Ƭvǁc�u�3���C���h�5���"�ӔҨ����7�w1 �Y�l�G��f�d���2�_ZT%7�=�UV���,'���hU��^�	fU��n�f�:��i ����#��a{[���i7�Cp�ؓb����y�D����s����=����"p8��ϱ����w/x�${�n����4j�	����Mhs��WZ���V�`�m����B#ڜF���F�D�h�Q��7B1�}N#Ɠ��V��~M��@ZO��,m�j���!_�!�d��艪�L}���"'��Mm��iB����s���p9Gz��;N]S����C[;�ɓ�F5�#�*�]�E�B���QʿK�$��"f�8.nG�<b�r��Wm����6�D�������B� ������������ոv9�?;��ͪ��T�/���М�s�;T:�Qg=&��Hb�>��F�?��������.��LE�\wf�#�'���:�&�O��b�6��P�S����x�0w�)Dx��Gr�0���u�Dw����F�Ĭ�Ns�>w�nz+����zL�%�\&*3�PyoA3b��)l�M�!a�HZ�V	ڵ��?��q���r�.��I�L�Z�k��+��F_av<�i7��d�	����l�G~��ѸFk�c�t���5�4G{�s�F&ְQ]��'��&��?#t�����N�����D�IWH��\��ҡ����_��I8wa:�P=mt�S�ik#L��n:��p��r�|>�.��>�5�F��ȉ��r"�VQ�DE9�y�?���[��J�ӑ+�VaF~�91מk�DlWvMG!�1sM�*���('D��v�B"�7T`�=��\����sw}���q�m��"Lim�֠�����C�3��j����K��#�!x��ĝ?b���ʱ�+�a�f�:\�G�Y��������*�Έ�;�/�,�d�>*�I��s'o�/��s�\C�3��;4�P(����������t̬(-��^V3����2��0}�[�px��{z��^�LwT��Dh��V������jUe��4O���Us��iJm���V�YJ�b(�{Uʣ�n����Y�\�vU�L�R{�W�x�n�<S)��<�<��[���l�dd�G�tx<��
����\>�\ꪬ���Ȓ��:٭8�DN��������rG�rx԰�N�2K=�5}��V���/��7�����cj�eU��*Y���J������;\N�Ȏ*���L9���,g���s���~��]�T����*�rF��y�&�=�^��iw;�urF�"�0y��.w�jd���B�v�|��1&_�e�V<>�W-��%{*�%��8S���"o�LΘ:)_�K��K���ty<��\���Q��^��%&�D���!S�Sz�.~���%��w�a�������n_��Q���v���V�'���ęy��jy��#W�dG��B��QJ�W�A�/p��>�s�Oq�aGq������u^�#۽�]�E=}�B��+����qxg	�(S����Z5�v7�=���%���*���U���*u9eQ�5 �,+�~�����U���e
Nh�����y���͔�vw��UE4�:S�s(�2M^��D��j�cm��rF�2��Ly��!n��:Q#.*���lq�}偃�ee��������v�������7��7?>��D�yq}3&M�]4��������NfVm�llL��6�q��7�B���eWs��k���Jf|y�)�~>H}7h~b����nF�aLJ�o~Jw��6�d�ym�&_uw�c��"M�Ƽ�y/�m��c1�h���E�7?jnI��k������0������I�&�H�e��/�u"�j�<)���QI��4���$��#Ѭ^|��o�7���/S�.�4�q��������~i�U.�U�O��ƉH�a��s.o3���E�z���z�HIy-V�<���Yy�!��Z�WD�9<���碖�Ga��o��~avO���k�a�D��0�ԯC��W��&~���&~��_"^����R��6��|�|�����7M5��"lh_6�}��Rp�<8�&'�mn��/��UٸX���/=|=�w��"~t��y����/��<�/���U����W��g"�_��~���&��"���`uC�މ�/�?������"~����W��#�����W�l�e���CE|&��E�j��S���<�_o�۴Q��i.
8���9�"��/ۮ�j|���?6 ަ���_�������E|���-%�z�J?uhX/�g��o��R����Us˧�J�S�����o��`��2M2�L�z��usK�?�z�M�]	R|�FɜoA���9�"MZ�}]�HkRDP3DZ|'Mv���
,3$Tw}�����n��yRb�I�,K��l'�Y�c6�5�2���u������2��t�H;/���SJ���W�Ep����M_�W��o�V?�c8(�.����\��z�h)׸Dl�r��q��y�罨"�lN姶I��6�±U�;�u�c,�����x��]yZ��_n�ь�$s�_���7�H�k�c�="��8v�F�/|b��s�%d>��dln�4h�(ʩA-�E�<)���Mʞ(e���/�2��,�&���SD�%�b���y��
E~>5�)���Ji�$�PJ-�6�y�YC���J�~1���"��8�D)�@�k�T���#��b�|�J�j�5Ζ�D@�?`���n_�V��ܒ�j��N��4�u�&Ѕ���;?�1Z�r-e�'H��V�6�"
stPa��1P��[�y�W�[��F;�z�/��Hs6;�]�7E���K�ˬ��ꑌ�6�y���c��f1V���]O6X�]x���GY��:\��(�?�?N�q�^�.;%��ժ�b�%����E��;Y�k�~ȇ�[��Ӥ��G��PP���S����b�꯰Ьo�Zb6�O1V��C"l�3L9�8�lX�~��"�������E��>[�Q_.�[�+��]�ǅ� �.�������fCO�3��8C���K��)�[���� ���7	�w�
�M���,�>�S�ב |���QB�.1��}R\��T�����:J��b�^}p��*��nl�����{���:� ~��$զ-(��W�҉g�c�=3�^7[�ĉcC�vv�3dwf����R��UI*�uP�j�P��R�ARE��Ҋ���Q��(�QZ��ʝ]�BԀ�?���K���~�>4�q�t���V,��0�xa�r����-���G��-[����k��T�y�Y]�nj�;Y~��Ѹ���^��3��䥛��R�8spԦ��4����lMٳ�0����Ap�֙~o��л�5[�������kF_ܺ�s^���f+��wm԰3}l>[͸���o��vp!˖���ݱ0̫ux��=xz۫[�k̶K�!���������`����|g�+��=����y��G����˷%�7��K������B?�u�4?X\t���j���,���0[�m/-ͮ_�FW�1��l�\����"������,?v�/���o�6�|C�n><��c[f������`y%(���>h7����]Z��W��\�{�h��'��ݧ��?��+���ť����`apo����/<����X��f7�m<�(^��_������Q8jܸn(^�������ʦ�sy�����/�?<��b�����Q;黮׾/�Ñ�Ƴ�5_}�����k�����/��|�[������͉���??5z7'ݱ��N��}�;��r՜8�'&[W5��a�8�p|<_�?lN�.�w������bo~y0tWJ��tW{�x�Zeb|���u����K��U�㍕��������hc�|�a6�:ꞱY�G,g���D�9��[�-dG���i�N�>�/8��؟�e���͉�p��6�;[��ya�;�;/�;/l�Fq����қ�-�z�������G{뜑�n,�6{+\���Ri��df��\6���wF��z`\�{|�����TltѸs�����^~$�K��:7Sֹ���L�9q�+�8��*I\-��|Rj'ݬT.��,ˢN�-?0��2ԥ�����J���ۥ�S��ѝ��,��a��0�֣��G�����a7L���Ds�RǕ�\�>_�T띸��Y�^�z�PyݚT��Zu�V-��R�è^�'ss�4ꔻ�N�Ӯm�d�_�J�uk�f�n�]	Ksݹ(?6YZʏTR��n')�+I�޾X����r7v��d�Jv��-i]����w �)���R��S�}��;��(�[>Q>Y�fyG孕J�ZiU�^���`�C��V>_��ʙ���a�
og�#ᯆO��~=<�3�+�Gǣ������蟣B|E���g�$�%����j�����?�g�-���O�K�I3�I$G��'�$�%M�~�Z�M�~����?��k�t*����������W�J����6��|�C�g�ۛ��w7כ��Z���í����ы�ѻ�=�w������������Wӗ�u]S��o��q�T�L������w�ᮟ��˻��~|�����{K�-����#�c�����t�K��4�h�h�͟n�|�Ps����懛_n�i���N��oE��ֻ[�����S��Z�n��o�<29;y��{&?0yr򣓟�ܼ��ޥ�Xy��L��*Q�r�|��!��3섽p�z�`�ះχ_�FWF�M��h-z(z$�����s�_G_��_?�e�W����/��ɭɡd6&����G��/&_I����\U}s�'�;�Q�U��������'�OU��~��7տ�~����k�kY���j��Gk/ԂtOz8���}����#��I�J?�>�~6�\���k�?����M�=}s}t^m�#ӰN���f�Ϳ�����R��5,����A������O��b """"""""""""""""""""""""""""""""�!{N<?v��oM�<]_?���}����u^��Ď��*�7xo��v|b���֯?��{f�~��Է�<2���=�gŇ���=SW�~z��w{��S[?޹m���ڱ+���P�r�����:��?v�������O_=uϓ/�͜������|>��������>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>������b�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|~�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�X���|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�_,��|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>��/�|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>���|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>����>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����������|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>������b�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|~�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�X���|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�_,��|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>��/�|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>���|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>����>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����������|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>������b�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|~�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����|>�����	   � ��E��~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������goH   qX��/����~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~���?{s@  �0���g~-������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~�ٛ   �A�?�h�~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������9   `�a�3�������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~����	   � ��E��~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������goH   qX��/����~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~���?{s@  �0���g~-������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~��������7$   �8�����~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������9   `�a�3�������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~����	   � ��E��~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������goH   qX��/����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~����  �a����"Z@������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~��������7$   �8�����~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������9   `�a�3�������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~����	   � ��E��~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~��������   0���_D����~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~����  �a����"Z@������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~��������7$   �8�����~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������9   `�a�3�������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~�ٛ   �A�?�h�~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~��������   0���_D����~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~����  �a����"Z@������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~��������7$   �8�����~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~���?{s@  �0���g~-������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~�ٛ   �A�?�h�~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~��������   0���_D����~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~����  �a����"Z@������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������goH   qX��/����~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~���?{s@  �0���g~-������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~�ٛ   �A�?�h�~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~��������   0���_D����~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~����	   � ��E��~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������goH   qX��/����~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~���?{s@  �0���g~-������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~�ٛ   �A�?�h�~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������9   `�a�3�������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~����	   � ��E��~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������goH   qX��/����~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~���?{s@  �0���g~-������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~��������7$   �8�����~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������9   `�a�3�������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~����	   � ��E��~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������goH   qX��/����~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~����  �a����"Z@������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~��������7$   �8�����~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������9   `�a�3�������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~����	   � ��E��~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~��������   0���_D����~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~����  �a����"Z@������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~��������7$   �8�����~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������9   `�a�3�������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�ٛ   �A�?�h�~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~��������   0���_D����~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~����  �a����"Z@������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~��������7$   �8�����~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���?{s@  �0���g~-������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~�ٛ   �A�?�h�~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~��������   0���_D����~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~����  �a����"Z@������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������goH   qX��/����~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~���?{s@  �0���g~-������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~�ٛ   �A�?�h�~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~��������   0���_D����~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����	   � ��E��~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������goH   qX��/����~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~���?{s@  �0���g~-������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~�ٛ   �A�?�h�~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������9   `�a�3������������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~����	   � ��E��~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������goH   qX��/����~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~���?{s@  �0���g~-������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~��������7$   �8�����~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������9   `�a�3�������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~����	   � ��E��~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������goH   qX��/����~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����  �a����"Z@���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~��������7$   �8�����~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������9   `�a�3�������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~����	   � ��E��~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~��������   0���_D���������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~����  �a����"Z@������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~��������7$   �8�����~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������9   `�a�3�������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�ٛ   �A�?�h������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~��������   0���_D����~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~����  �a����"Z@������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~��������7$   �8�����~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���?{s@  �0���g~-����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~�ٛ   �A�?�h�~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~��������   0���_D����~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~����  �a����"Z@������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������goH   qX��/�l~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~���?{s@  �0���g~-������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~�ٛ   �A�?�h�~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~��������   0���_D����~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~goH   1x��/������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�߿�~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����/������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�߿�~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����/������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�߿�~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����/������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�߿�~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����/������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�߿�~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����/������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�߿�~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����/������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�߿�~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����/������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�߿�~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����/������~������~������~������~������~������~������~������~������~������~������~��������7$   �8�����~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������9   `�a�3�������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~����	   � ��E��~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���ogoH   qX��/����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~����  �a����"Z@������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~��������7$   �8�����~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������9   `�a�3�������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���������	   � ��E��~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~��������   0���_D����~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~����  �a����"Z@������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~��������7$   �8�����~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������9   `�a�3�������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~�ٛ   �A�?�h�~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~��������   0���_D����~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~����  �a����"Z@������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������7$   �8�����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~���?{s@  �0���g~-������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~�ٛ   �A�?�h�~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~��������   0���_D����~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~����  �a����"Z@������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������goH   qX��/����~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~���?{s@  �0���g~-������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~�ٛ   �A�?�h�~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�������������   0���_D����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~����	   � ��E��~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������goH   qX��/����~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~���?{s@  �0���g~-������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~�ٛ   �A�?�h�~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������9   `�a�3�������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~����	   � ��E��~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������goH   qX��/����~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~���?{s@  �0���g~-������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~��������7$   �8�����~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������9   `�a�3�������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~����	   � ��E��~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������goH   qX��/����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~����  �a����"Z@������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~��������7$   �8�����~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������9   `�a�3�������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~����	   � ��E��~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~��������   0���_D����~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~����  �a����"Z@������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~��������7$   �8�����~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������9   `�a�3�������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~�ٛ   �A�?�h�~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~��������   0���_D����~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~����  �a����"Z@������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~��������7$   �8�����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~���?{s@  �0���g~-������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~�ٛ   �A�?�h�~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~��������   0���_D����~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~����  �a����"Z@������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������goH   qX��/����~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~���?{s@  �0���g~-������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~�ٛ   �A�?�h�~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~��������   0���_D����~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~����	   � ��E��~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������goH   qX��/����~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~���?{s@  �0���g~-������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~�ٛ   �A�?�h�~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������9   `�a�3�������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~����	   � ��E��~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������goH   qX��/����~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~���?{s@  �0���g~-������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~��������7$   �8�����~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������9   `�a�3�������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~����	   � ��E��~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������goH   qX��/����~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~����  �a����"Z@������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~��������7$   �8�����~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������9   `�a�3�������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~����	   � ��E��~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~��������   0���_D����~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~����  �a����"Z@������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~��������7$   �8�����~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������9   `�a�3�������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�ٛ   �A�?�h�~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~��������   0���_D����~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~����  �a����"Z@������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~��������7$   �8�����~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~���?{s@  �0���g~-������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~�ٛ   �A�?�h�~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~��������   0���_D����~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~����  �a����"Z@������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������goH   qX��/����~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~���?{s@  �0���g~-������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~�ٛ   �A�?�h�~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~��������   0���_D����~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����	   � ��E��~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������goH   qX��/����~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~���?{s@  �0���g~-������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~�ٛ   �A�?�h�~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������9   `�a�3�������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~����	   � ��E��~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������goH   qX��/����~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~���?{s@  �0���g~-������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~��������7$   �8�����~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������9   `�a�3�������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~����	   � ��E��~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������goH   qX��/����~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����  �a����"Z@�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~��������7$   �8�����~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������9   `�a�3�������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~����	   � ��E��~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~��������   0���_D���������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~����  �a����"Z@������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~��������7$   �8�����~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������9   `�a�3�������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�ٛ   �A�?�h�~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~��������   0���_D����~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~����  �a����"Z@������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~��������7$   �8�����~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���?{s@  �0���g~-���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~�ٛ   �A�?�h�~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~��������   0���_D����~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~����  �a����"Z@������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������goH   qX��/���������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~���?{s@  �0���g~-������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~�ٛ   �A�?�h�~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~��������   0���_D����~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����	   � ��E�������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������goH   qX��/����~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~���?{s@  �0���g~-������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~�ٛ   �A�?�h�~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������9   `�a�3�����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~����	   � ��E��~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������goH   qX��/����~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~���?{s@  �0���g~-������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~��������9   `���3��0������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�߿�~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����/������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�߿�~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����/������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�߿�~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����/������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�߿�~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����/������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�߿�~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����/������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�߿�~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����/������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�߿�~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����/������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�߿�~������~������~������~������~������~������~������~������~������~������~������~��������   0���_D����~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~����  �a����"Z@������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~��������7$   �8�����~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����9   `�a�3�������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~�ٛ   �A�?�h�~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~��������   0���_D����~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~����  �a����"Z@������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o��7$   �8�����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~���?{s@  �0���g~-������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~�ٛ   �A�?�h�~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~��������   0���_D����~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���������  �a����"Z@������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������goH   qX��/����~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~���?{s@  �0���g~-������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~�ٛ   �A�?�h�~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�������������   0���_D����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~����	   � ��E��~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������goH   qX��/����~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~���?{s@  �0���g~-������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~�ٛ   �A�?�h�~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������9   `�a�3�������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~����	   � ��E��~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������goH   qX��/����~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~���?{s@  �0���g~-������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~��������7$   �8�����~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������9   `�a�3�������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~����	   � ��E��~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������goH   qX��/����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~����  �a����"Z@������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~��������7$   �8�����~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������9   `�a�3�������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~����	   � ��E��~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~��������   0���_D����~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~����  �a����"Z@������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~��������7$   �8�����~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������9   `�a�3�������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~�ٛ   �A�?�h�~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~��������   0���_D����~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~����  �a����"Z@������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~��������7$   �8�����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~���?{s@  �0���g~-������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~�ٛ   �A�?�h�~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~��������   0���_D����~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~����  �a����"Z@������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������goH   qX��/����~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~���?{s@  �0���g~-������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~�ٛ   �A�?�h�~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~��������   0���_D����~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~����	   � ��E��~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������goH   qX��/����~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~���?{s@  �0���g~-������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~�ٛ   �A�?�h�~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������9   `�a�3�������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~����	   � ��E��~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������goH   qX��/����~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~���?{s@  �0���g~-������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~��������7$   �8�����~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������9   `�a�3�������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~����	   � ��E��~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������goH   qX��/����~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~����  �a����"Z@������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~��������7$   �8�����~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������9   `�a�3�������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~����	   � ��E��~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~��������   0���_D����~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~����  �a����"Z@������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~��������7$   �8�����~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������9   `�a�3�������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~�ٛ   �A�?�h�~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~��������   0���_D����~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~����  �a����"Z@������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~��������7$   �8�����~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~���?{s@  �0���g~-������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~�ٛ   �A�?�h�~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~��������   0���_D����~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~����  �a����"Z@������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������goH   qX��/����~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~���?{s@  �0���g~-������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~�ٛ   �A�?�h�~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~��������   0���_D����~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����	   � ��E��~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������goH   qX��/����~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~���?{s@  �0���g~-������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~�ٛ   �A�?�h�~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������9   `�a�3�������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~����	   � ��E��~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������goH   qX��/����~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~���?{s@  �0���g~-������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~��������7$   �8�����~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������9   `�a�3�������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~����	   � ��E��~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������goH   qX��/����~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����  �a����"Z@�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~��������7$   �8�����~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������9   `�a�3�������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~����	   � ��E��~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~��������   0���_D����~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~����  �a����"Z@������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~��������7$   �8�����~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������9   `�a�3�������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�ٛ   �A�?�h�~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~��������   0���_D����~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~����  �a����"Z@������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~��������7$   �8�����~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���?{s@  �0���g~-�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~�ٛ   �A�?�h�~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~��������   0���_D����~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~����  �a����"Z@������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������goH   qX��/���������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~���?{s@  �0���g~-������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~�ٛ   �A�?�h�~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~��������   0���_D����~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����	   � ��E��~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������goH   qX��/����~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~���?{s@  �0���g~-������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~�ٛ   �A�?�h�~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������9   `�a�3����o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~����	   � ��E��~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������goH   qX��/����~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~���?{s@  �0���g~-������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~��������7$   �8����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������9   `�a�3�������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~����	   � ��E��~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������goH   qX��/����~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����  �a����"Z�����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~��������7$   �8�����~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������9   `�a�3�������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~����	   � ��E��~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����w��  �a����"Z��~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����/������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�߿�~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����/������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�߿�~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����/������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�߿�~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����/������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�߿�~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����/������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�߿�~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����/������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�߿�~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����/������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�߿�~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����/������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~���?{s@  �0���g~-������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~�ٛ   �A�?�h�~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~��������   0���_D����~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�������v��  �a����"Z@������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������goH   qX��/����~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~���?{s@  �0���g~-������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~�ٛ   �A�?�h�~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������   0���_D����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~����	   � ��E��~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������goH   qX��/����~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~���?{s@  �0���g~-������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~�ٛ   �A�?�h�~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������9   `�a�3�������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~����	   � ��E��~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������goH   qX��/����~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~��������?{s@  �0���g~-������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~��������7$   �8�����~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������9   `�a�3�������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~����	   � ��E��~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������goH   qX��/����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~����  �a����"Z@������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~��������7$   �8�����~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������9   `�a�3�������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~����	   � ��E��~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~��������   0���_D����~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~����  �a����"Z@������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~��������7$   �8�����~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������9   `�a�3�������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~�ٛ   �A�?�h�~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~��������   0���_D����~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~����  �a����"Z@������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�������������7$   �8�����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~���?{s@  �0���g~-������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~�ٛ   �A�?�h�~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~��������   0���_D����~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~����  �a����"Z@������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������goH   qX��/����~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~���?{s@  �0���g~-������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~�ٛ   �A�?�h�~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~��������   0���_D����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~����	   � ��E��~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������goH   qX��/����~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~���?{s@  �0���g~-������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~�ٛ   �A�?�h�~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������9   `�a�3�������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~����	   � ��E��~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������goH   qX��/����~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~���?{s@  �0���g~-������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~��������7$   �8�����~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������9   `�a�3�������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~����	   � ��E��~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������goH   qX��/����~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~����  �a����"Z@������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~��������7$   �8�����~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������9   `�a�3�������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~����	   � ��E��~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~��������   0���_D����~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~����  �a����"Z@������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~��������7$   �8�����~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������9   `�a�3�������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~�ٛ   �A�?�h�~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~��������   0���_D����~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~����  �a����"Z@������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~��������7$   �8�����~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~���?{s@  �0���g~-������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~�ٛ   �A�?�h�~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~��������   0���_D����~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~����  �a����"Z@������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������goH   qX��/����~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~���?{s@  �0���g~-������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~�ٛ   �A�?�h�~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~��������   0���_D����~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~����	   � ��E��~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������goH   qX��/����~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~���?{s@  �0���g~-������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~�ٛ   �A�?�h�~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������9   `�a�3�������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~����	   � ��E��~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������goH   qX��/����~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~���?{s@  �0���g~-������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~��������7$   �8�����~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������9   `�a�3�������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~����	   � ��E��~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������goH   qX��/����~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����  �a����"Z@������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~��������7$   �8�����~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������9   `�a�3�������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~����	   � ��E��~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~��������   0���_D����~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~����  �a����"Z@������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~��������7$   �8�����~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������9   `�a�3�������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�ٛ   �A�?�h�~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~��������   0���_D����~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~����  �a����"Z@������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~��������7$   �8�����~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���?{s@  �0���g~-�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~�ٛ   �A�?�h�~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~��������   0���_D����~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~����  �a����"Z@������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������goH   qX��/����~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~���?{s@  �0���g~-������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~�ٛ   �A�?�h�~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~��������   0���_D����~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����	   � ��E��~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������goH   qX��/����~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~���?{s@  �0���g~-������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~�ٛ   �A�?�h�~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������9   `�a�3������������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~����	   � ��E��~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������goH   qX��/����~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~���?{s@  �0���g~-������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~��������7$   �8����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������9   `�a�3�������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~����	   � ��E��~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������goH   qX��/����~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����  �a����"Z@����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~��������7$   �8�����~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������9   `�a�3�������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~����	   � ��E��~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~��������   0���_D�o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~����  �a����"Z@������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~��������7$   �8�����~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������9   `�a�3�������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�ٛ   �A�?�h������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~��������   0���_D����~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~����  �a����"Z@������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~��������7$   �8�����~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���ٛ   �A�?�h���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�߿�~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����/������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�߿�~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����/������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�߿�~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����/������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�߿�~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����/������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�߿�~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����/������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�߿�~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����/������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�߿�~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����/������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�߿�~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����/������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~����	   � ��E��~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������goH   qX��/����~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~���?{s@  �0���g~-������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������ٛ   �A�?�h�~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������9   `�a�3�������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~����	   � ��E��~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������goH   qX��/����~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~��������?{s@  �0���g~-������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~��������7$   �8�����~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������9   `�a�3�������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~����	   � ��E��~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����goH   qX��/����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~����  �a����"Z@������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~��������7$   �8�����~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������9   `�a�3�������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~����	   � ��E��~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~��������   0���_D����~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~����  �a����"Z@������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~��������7$   �8�����~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������9   `�a�3�������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~�ٛ   �A�?�h�~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~��������   0���_D����~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~����  �a����"Z@������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�������������7$   �8�����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~���?{s@  �0���g~-������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~�ٛ   �A�?�h�~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~��������   0���_D����~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~����  �a����"Z@������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������goH   qX��/����~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~���?{s@  �0���g~-������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~�ٛ   �A�?�h�~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~��������   0���_D����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~����	   � ��E��~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������goH   qX��/����~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~���?{s@  �0���g~-������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~�ٛ   �A�?�h�~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������9   `�a�3�������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~����	   � ��E��~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������goH   qX��/����~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~���?{s@  �0���g~-������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~��������7$   �8�����~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������9   `�a�3�������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~����	   � ��E��~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������goH   qX��/����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~����  �a����"Z@������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~��������7$   �8�����~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������9   `�a�3�������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~����	   � ��E��~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~��������   0���_D����~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~����  �a����"Z@������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~��������7$   �8�����~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������9   `�a�3�������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~�ٛ   �A�?�h�~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~��������   0���_D����~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~����  �a����"Z@������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~��������7$   �8�����~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~���?{s@  �0���g~-������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~�ٛ   �A�?�h�~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~��������   0���_D����~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~����  �a����"Z@������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������goH   qX��/����~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~���?{s@  �0���g~-������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~�ٛ   �A�?�h�~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~��������   0���_D����~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~����	   � ��E��~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������goH   qX��/����~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~���?{s@  �0���g~-������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~�ٛ   �A�?�h�~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������9   `�a�3�������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~����	   � ��E��~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������goH   qX��/����~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~���?{s@  �0���g~-������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~��������7$   �8�����~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������9   `�a�3�������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~����	   � ��E��~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������goH   qX��/����~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~����  �a����"Z@������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~��������7$   �8�����~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������9   `�a�3�������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~����	   � ��E��~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~��������   0���_D����~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~����  �a����"Z@������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~��������7$   �8�����~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������9   `�a�3�������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�ٛ   �A�?�h�~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~��������   0���_D����~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~����  �a����"Z@������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~��������7$   �8�����~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���?{s@  �0���g~-������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~�ٛ   �A�?�h�~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~��������   0���_D����~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~����  �a����"Z@������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������goH   qX��/����~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~���?{s@  �0���g~-������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~�ٛ   �A�?�h�~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~��������   0���_D����~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����	   � ��E��~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������goH   qX��/����~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~���?{s@  �0���g~-������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~�ٛ   �A�?�h�~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������9   `�a�3������������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~����	   � ��E��~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������goH   qX��/����~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~���?{s@  �0���g~-������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~��������7$   �8�����~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������9   `�a�3�������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~����	   � ��E��~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������goH   qX��/����~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����  �a����"Z@���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~��������7$   �8�����~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������9   `�a�3�������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~����	   � ��E��~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~��������   0���_D���������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~����  �a����"Z@������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~��������7$   �8�����~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������9   `�a�3�������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�ٛ   �A�?�h������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~��������   0���_D����~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~����  �a����"Z@������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~��������7$   �8�����~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���?{s@  �0���g~-����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~�ٛ   �A�?�h�~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~��������   0���_D����~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~����  �a����"Z@������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������goH   qX��/�l~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~���?{s@  �0���g~-������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~�ٛ   �A�?�h�~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~��������   0���_D����~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~goH   1x��/������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�߿�~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����/������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�߿�~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����/������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�߿�~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����/������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�߿�~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����/������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�߿�~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����/������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�߿�~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����/������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�߿�~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����/������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�߿�~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����/������~������~������~������~������~������~������~������~������~������~������~��������7$   �8�����~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������9   `�a�3�������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~����	   � ��E��~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���ogoH   qX��/����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~����  �a����"Z@������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~��������7$   �8�����~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������9   `�a�3�������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���������	   � ��E��~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~��������   0���_D����~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~����  �a����"Z@������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~��������7$   �8�����~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������9   `�a�3�������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~�ٛ   �A�?�h�~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~��������   0���_D����~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~����  �a����"Z@������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������7$   �8�����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~���?{s@  �0���g~-������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~�ٛ   �A�?�h�~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~��������   0���_D����~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~����  �a����"Z@������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������goH   qX��/����~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~���?{s@  �0���g~-������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~�ٛ   �A�?�h�~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�������������   0���_D����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~����	   � ��E��~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������goH   qX��/����~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~���?{s@  �0���g~-������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~�ٛ   �A�?�h�~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������9   `�a�3�������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~����	   � ��E��~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������goH   qX��/����~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~���?{s@  �0���g~-������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~��������7$   �8�����~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������9   `�a�3�������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~����	   � ��E��~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������goH   qX��/����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~����  �a����"Z@������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~��������7$   �8�����~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������9   `�a�3�������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~����	   � ��E��~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~��������   0���_D����~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~����  �a����"Z@������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~��������7$   �8�����~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������9   `�a�3�������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~�ٛ   �A�?�h�~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~��������   0���_D����~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~����  �a����"Z@������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~��������7$   �8�����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~���?{s@  �0���g~-������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~�ٛ   �A�?�h�~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~��������   0���_D����~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~����  �a����"Z@������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������goH   qX��/����~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~���?{s@  �0���g~-������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~�ٛ   �A�?�h�~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~��������   0���_D����~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~����	   � ��E��~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������goH   qX��/����~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~���?{s@  �0���g~-������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~�ٛ   �A�?�h�~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������9   `�a�3�������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~����	   � ��E��~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������goH   qX��/����~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~���?{s@  �0���g~-������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~��������7$   �8�����~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������9   `�a�3�������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~����	   � ��E��~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������goH   qX��/����~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~����  �a����"Z@������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~��������7$   �8�����~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������9   `�a�3�������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~����	   � ��E��~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~��������   0���_D����~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~����  �a����"Z@������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~��������7$   �8�����~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������9   `�a�3�������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�ٛ   �A�?�h�~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~��������   0���_D����~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~����  �a����"Z@������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~��������7$   �8�����~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~���?{s@  �0���g~-������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~�ٛ   �A�?�h�~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~��������   0���_D����~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~����  �a����"Z@������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������goH   qX��/����~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~���?{s@  �0���g~-������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~�ٛ   �A�?�h�~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~��������   0���_D����~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����	   � ��E��~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������goH   qX��/����~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~���?{s@  �0���g~-������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~�ٛ   �A�?�h�~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������9   `�a�3�������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~����	   � ��E��~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������goH   qX��/����~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~���?{s@  �0���g~-������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~��������7$   �8�����~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������9   `�a�3�������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~����	   � ��E��~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������goH   qX��/����~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����  �a����"Z@�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~��������7$   �8�����~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������9   `�a�3�������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~����	   � ��E��~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~��������   0���_D���������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~����  �a����"Z@������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~��������7$   �8�����~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������9   `�a�3�������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�ٛ   �A�?�h�~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~��������   0���_D����~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~����  �a����"Z@������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~��������7$   �8�����~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���?{s@  �0���g~-���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~�ٛ   �A�?�h�~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~��������   0���_D����~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~����  �a����"Z@������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������goH   qX��/���������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~���?{s@  �0���g~-������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~�ٛ   �A�?�h�~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~��������   0���_D����~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����	   � ��E�������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������goH   qX��/����~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~���?{s@  �0���g~-������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~�ٛ   �A�?�h�~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������9   `�a�3�����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~����	   � ��E��~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������goH   qX��/����~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~���?{s@  �0���g~-������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~��������9   `���3��0������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�߿�~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����/������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�߿�~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����/������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�߿�~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����/������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�߿�~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����/������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�߿�~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����/������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�߿�~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����/������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�߿�~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����/������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�߿�~������~������~������~������~������~������~������~������~������~������~������~��������   0���_D����~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~����  �a����"Z@������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~��������7$   �8�����~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����9   `�a�3�������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~�ٛ   �A�?�h�~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~��������   0���_D����~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~����  �a����"Z@������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o��7$   �8�����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~���?{s@  �0���g~-������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~�ٛ   �A�?�h�~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~��������   0���_D����~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���������  �a����"Z@������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������goH   qX��/����~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~���?{s@  �0���g~-������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~�ٛ   �A�?�h�~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�������������   0���_D����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~����	   � ��E��~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������goH   qX��/����~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~���?{s@  �0���g~-������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~�ٛ   �A�?�h�~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������9   `�a�3�������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~����	   � ��E��~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������goH   qX��/����~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~���?{s@  �0���g~-������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~��������7$   �8�����~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������9   `�a�3�������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~����	   � ��E��~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������goH   qX��/����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~����  �a����"Z@������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~��������7$   �8�����~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������9   `�a�3�������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~����	   � ��E��~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~��������   0���_D����~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~����  �a����"Z@������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~��������7$   �8�����~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������9   `�a�3�������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~�ٛ   �A�?�h�~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~��������   0���_D����~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~����  �a����"Z@������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~��������7$   �8�����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~���?{s@  �0���g~-������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~�ٛ   �A�?�h�~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~��������   0���_D����~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~����  �a����"Z@������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������goH   qX��/����~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~���?{s@  �0���g~-������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~�ٛ   �A�?�h�~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~��������   0���_D����~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~����	   � ��E��~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������goH   qX��/����~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~���?{s@  �0���g~-������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~�ٛ   �A�?�h�~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������9   `�a�3�������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~����	   � ��E��~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������goH   qX��/����~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~���?{s@  �0���g~-������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~��������7$   �8�����~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������9   `�a�3�������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~����	   � ��E��~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������goH   qX��/����~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~����  �a����"Z@������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~��������7$   �8�����~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������9   `�a�3�������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~����	   � ��E��~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~��������   0���_D����~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~����  �a����"Z@������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~��������7$   �8�����~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������9   `�a�3�������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~�ٛ   �A�?�h�~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~��������   0���_D����~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~����  �a����"Z@������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~��������7$   �8�����~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~���?{s@  �0���g~-������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~�ٛ   �A�?�h�~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~��������   0���_D����~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~����  �a����"Z@������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������goH   qX��/����~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~���?{s@  �0���g~-������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~�ٛ   �A�?�h�~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~��������   0���_D����~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����	   � ��E��~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������goH   qX��/����~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~���?{s@  �0���g~-������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~�ٛ   �A�?�h�~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������9   `�a�3�������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~����	   � ��E��~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������goH   qX��/����~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~���?{s@  �0���g~-������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~��������7$   �8�����~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������9   `�a�3�������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~����	   � ��E��~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������goH   qX��/����~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����  �a����"Z@�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~��������7$   �8�����~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������9   `�a�3�������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~����	   � ��E��~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~��������   0���_D����~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~����  �a����"Z@������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~��������7$   �8�����~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������9   `�a�3�������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�ٛ   �A�?�h�~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~��������   0���_D����~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~����  �a����"Z@������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~��������7$   �8�����~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���?{s@  �0���g~-�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~�ٛ   �A�?�h�~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~��������   0���_D����~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~����  �a����"Z@������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������goH   qX��/���������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~���?{s@  �0���g~-������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~�ٛ   �A�?�h�~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~��������   0���_D����~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����	   � ��E��~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������goH   qX��/����~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~���?{s@  �0���g~-������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~�ٛ   �A�?�h�~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������9   `�a�3����o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~����	   � ��E��~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������goH   qX��/����~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~���?{s@  �0���g~-������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~��������7$   �8����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������9   `�a�3�������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~����	   � ��E��~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������goH   qX��/����~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����  �a����"Z�����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~��������7$   �8�����~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������9   `�a�3�������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~����	   � ��E��~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����w��  �a����"Z��~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����/������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�߿�~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����/������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�߿�~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����/������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�߿�~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����/������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�߿�~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����/������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�߿�~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����/������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�߿�~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����/������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�߿�~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����/������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~���?{s@  �0���g~-������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~�ٛ   �A�?�h�~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~��������   0���_D����~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�������v��  �a����"Z@������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������goH   qX��/����~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~���?{s@  �0���g~-������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~�ٛ   �A�?�h�~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������   0���_D����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~����	   � ��E��~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������goH   qX��/����~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~���?{s@  �0���g~-������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~�ٛ   �A�?�h�~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������9   `�a�3�������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~����	   � ��E��~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������goH   qX��/����~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~��������?{s@  �0���g~-������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~��������7$   �8�����~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������9   `�a�3�������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~����	   � ��E��~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������goH   qX��/����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~����  �a����"Z@������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~��������7$   �8�����~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������9   `�a�3�������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~����	   � ��E��~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~��������   0���_D����~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~����  �a����"Z@������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~��������7$   �8�����~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������9   `�a�3�������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~�ٛ   �A�?�h�~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~��������   0���_D����~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~����  �a����"Z@������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�������������7$   �8�����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~���?{s@  �0���g~-������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~�ٛ   �A�?�h�~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~��������   0���_D����~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~����  �a����"Z@������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������goH   qX��/����~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~���?{s@  �0���g~-������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~�ٛ   �A�?�h�~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~��������   0���_D����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~����	   � ��E��~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������goH   qX��/����~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~���?{s@  �0���g~-������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~�ٛ   �A�?�h�~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������9   `�a�3�������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~����	   � ��E��~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������goH   qX��/����~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~���?{s@  �0���g~-������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~��������7$   �8�����~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������9   `�a�3�������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~����	   � ��E��~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������goH   qX��/����~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~����  �a����"Z@������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~��������7$   �8�����~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������9   `�a�3�������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~����	   � ��E��~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~��������   0���_D����~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~����  �a����"Z@������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~��������7$   �8�����~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������9   `�a�3�������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~�ٛ   �A�?�h�~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~��������   0���_D����~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~����  �a����"Z@������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~��������7$   �8�����~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~���?{s@  �0���g~-������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~�ٛ   �A�?�h�~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~��������   0���_D����~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~����  �a����"Z@������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������goH   qX��/����~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~���?{s@  �0���g~-������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~�ٛ   �A�?�h�~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~��������   0���_D����~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~����	   � ��E��~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������goH   qX��/����~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~���?{s@  �0���g~-������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~�ٛ   �A�?�h�~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������9   `�a�3�������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~����	   � ��E��~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������goH   qX��/����~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~���?{s@  �0���g~-������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~��������7$   �8�����~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������9   `�a�3�������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~����	   � ��E��~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������goH   qX��/����~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����  �a����"Z@������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~��������7$   �8�����~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������9   `�a�3�������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~����	   � ��E��~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~��������   0���_D����~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~����  �a����"Z@������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~��������7$   �8�����~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������9   `�a�3�������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�ٛ   �A�?�h�~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~��������   0���_D����~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~����  �a����"Z@������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~��������7$   �8�����~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���?{s@  �0���g~-�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~�ٛ   �A�?�h�~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~��������   0���_D����~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~����  �a����"Z@������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������goH   qX��/����~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~���?{s@  �0���g~-������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~�ٛ   �A�?�h�~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~��������   0���_D����~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����	   � ��E��~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������goH   qX��/����~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~���?{s@  �0���g~-������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~�ٛ   �A�?�h�~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������9   `�a�3������������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~����	   � ��E��~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������goH   qX��/����~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~���?{s@  �0���g~-������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����7������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���~������~������~������~������~������~������~������~������~������~������~������~������~������~������~��������75  0����k��=� ~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~���o~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~�����������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~������~����~������~������~������~������~������~�������~������~������~������~������~��������������~������~������~������~������~�������~������~������~������~������~������~�������~������~������~������~������~������~�������~������~������~������~������~��������������~������~������~������~������~�������~������~������~������~������~������~�����PK 
     !F�V             $              new/
         ����ފ���}�ފ�����ފ�PK     ���Ve��2�6 �o= $           "   new/SETUP.exe
         �,Y-���w��ފ�w��ފ�PK      �   �6   